// Stub master driver BFM - replace with actual implementation
interface axi4_master_driver_bfm(input aclk, input aresetn);
endinterface
