// Stub slave driver BFM - replace with actual implementation
interface axi4_slave_driver_bfm(input aclk, input aresetn);
endinterface
