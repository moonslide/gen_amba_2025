// Stub master monitor BFM - replace with actual implementation
module axi4_master_monitor_bfm(input aclk, input aresetn);
endmodule
