//==============================================================================
// axi4_master_seq_pkg.sv
// Generated for 16x16 VIP RTL Integration
// Date: 2025-08-06 22:49:41
//==============================================================================

package axi4_master_seq_pkg;
    
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import axi4_globals_pkg::*;
    import axi4_master_pkg::*;
    
    // Include all sequence files
    `include "axi4_master_base_seq.sv"
    `include "axi4_master_write_seq.sv"
    `include "axi4_master_read_seq.sv"
    `include "axi4_master_burst_seq.sv"
    `include "axi4_master_random_seq.sv"
    `include "axi4_master_qos_seq.sv"
    
endpackage : axi4_master_seq_pkg
