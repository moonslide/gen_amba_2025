// Master 1 connections
,.m1_awid(rtl_m_awid[1]), .m1_awaddr(rtl_m_awaddr[1]), .m1_awlen(rtl_m_awlen[1]),
.m1_awsize(rtl_m_awsize[1]), .m1_awburst(rtl_m_awburst[1]), .m1_awlock(rtl_m_awlock[1]),
.m1_awcache(rtl_m_awcache[1]), .m1_awprot(rtl_m_awprot[1]), .m1_awqos(rtl_m_awqos[1]),
.m1_awvalid(rtl_m_awvalid[1]), .m1_awready(rtl_m_awready[1]),
.m1_wdata(rtl_m_wdata[1]), .m1_wstrb(rtl_m_wstrb[1]), .m1_wlast(rtl_m_wlast[1]),
.m1_wvalid(rtl_m_wvalid[1]), .m1_wready(rtl_m_wready[1]),
.m1_bid(rtl_m_bid[1]), .m1_bresp(rtl_m_bresp[1]), .m1_bvalid(rtl_m_bvalid[1]), .m1_bready(rtl_m_bready[1]),
.m1_arid(rtl_m_arid[1]), .m1_araddr(rtl_m_araddr[1]), .m1_arlen(rtl_m_arlen[1]),
.m1_arsize(rtl_m_arsize[1]), .m1_arburst(rtl_m_arburst[1]), .m1_arlock(rtl_m_arlock[1]),
.m1_arcache(rtl_m_arcache[1]), .m1_arprot(rtl_m_arprot[1]), .m1_arqos(rtl_m_arqos[1]),
.m1_arvalid(rtl_m_arvalid[1]), .m1_arready(rtl_m_arready[1]),
.m1_rid(rtl_m_rid[1]), .m1_rdata(rtl_m_rdata[1]), .m1_rresp(rtl_m_rresp[1]),
.m1_rlast(rtl_m_rlast[1]), .m1_rvalid(rtl_m_rvalid[1]), .m1_rready(rtl_m_rready[1]),

// Master 2 connections
.m2_awid(rtl_m_awid[2]), .m2_awaddr(rtl_m_awaddr[2]), .m2_awlen(rtl_m_awlen[2]),
.m2_awsize(rtl_m_awsize[2]), .m2_awburst(rtl_m_awburst[2]), .m2_awlock(rtl_m_awlock[2]),
.m2_awcache(rtl_m_awcache[2]), .m2_awprot(rtl_m_awprot[2]), .m2_awqos(rtl_m_awqos[2]),
.m2_awvalid(rtl_m_awvalid[2]), .m2_awready(rtl_m_awready[2]),
.m2_wdata(rtl_m_wdata[2]), .m2_wstrb(rtl_m_wstrb[2]), .m2_wlast(rtl_m_wlast[2]),
.m2_wvalid(rtl_m_wvalid[2]), .m2_wready(rtl_m_wready[2]),
.m2_bid(rtl_m_bid[2]), .m2_bresp(rtl_m_bresp[2]), .m2_bvalid(rtl_m_bvalid[2]), .m2_bready(rtl_m_bready[2]),
.m2_arid(rtl_m_arid[2]), .m2_araddr(rtl_m_araddr[2]), .m2_arlen(rtl_m_arlen[2]),
.m2_arsize(rtl_m_arsize[2]), .m2_arburst(rtl_m_arburst[2]), .m2_arlock(rtl_m_arlock[2]),
.m2_arcache(rtl_m_arcache[2]), .m2_arprot(rtl_m_arprot[2]), .m2_arqos(rtl_m_arqos[2]),
.m2_arvalid(rtl_m_arvalid[2]), .m2_arready(rtl_m_arready[2]),
.m2_rid(rtl_m_rid[2]), .m2_rdata(rtl_m_rdata[2]), .m2_rresp(rtl_m_rresp[2]),
.m2_rlast(rtl_m_rlast[2]), .m2_rvalid(rtl_m_rvalid[2]), .m2_rready(rtl_m_rready[2]),

// Master 3 connections
.m3_awid(rtl_m_awid[3]), .m3_awaddr(rtl_m_awaddr[3]), .m3_awlen(rtl_m_awlen[3]),
.m3_awsize(rtl_m_awsize[3]), .m3_awburst(rtl_m_awburst[3]), .m3_awlock(rtl_m_awlock[3]),
.m3_awcache(rtl_m_awcache[3]), .m3_awprot(rtl_m_awprot[3]), .m3_awqos(rtl_m_awqos[3]),
.m3_awvalid(rtl_m_awvalid[3]), .m3_awready(rtl_m_awready[3]),
.m3_wdata(rtl_m_wdata[3]), .m3_wstrb(rtl_m_wstrb[3]), .m3_wlast(rtl_m_wlast[3]),
.m3_wvalid(rtl_m_wvalid[3]), .m3_wready(rtl_m_wready[3]),
.m3_bid(rtl_m_bid[3]), .m3_bresp(rtl_m_bresp[3]), .m3_bvalid(rtl_m_bvalid[3]), .m3_bready(rtl_m_bready[3]),
.m3_arid(rtl_m_arid[3]), .m3_araddr(rtl_m_araddr[3]), .m3_arlen(rtl_m_arlen[3]),
.m3_arsize(rtl_m_arsize[3]), .m3_arburst(rtl_m_arburst[3]), .m3_arlock(rtl_m_arlock[3]),
.m3_arcache(rtl_m_arcache[3]), .m3_arprot(rtl_m_arprot[3]), .m3_arqos(rtl_m_arqos[3]),
.m3_arvalid(rtl_m_arvalid[3]), .m3_arready(rtl_m_arready[3]),
.m3_rid(rtl_m_rid[3]), .m3_rdata(rtl_m_rdata[3]), .m3_rresp(rtl_m_rresp[3]),
.m3_rlast(rtl_m_rlast[3]), .m3_rvalid(rtl_m_rvalid[3]), .m3_rready(rtl_m_rready[3]),

// Master 4 connections
.m4_awid(rtl_m_awid[4]), .m4_awaddr(rtl_m_awaddr[4]), .m4_awlen(rtl_m_awlen[4]),
.m4_awsize(rtl_m_awsize[4]), .m4_awburst(rtl_m_awburst[4]), .m4_awlock(rtl_m_awlock[4]),
.m4_awcache(rtl_m_awcache[4]), .m4_awprot(rtl_m_awprot[4]), .m4_awqos(rtl_m_awqos[4]),
.m4_awvalid(rtl_m_awvalid[4]), .m4_awready(rtl_m_awready[4]),
.m4_wdata(rtl_m_wdata[4]), .m4_wstrb(rtl_m_wstrb[4]), .m4_wlast(rtl_m_wlast[4]),
.m4_wvalid(rtl_m_wvalid[4]), .m4_wready(rtl_m_wready[4]),
.m4_bid(rtl_m_bid[4]), .m4_bresp(rtl_m_bresp[4]), .m4_bvalid(rtl_m_bvalid[4]), .m4_bready(rtl_m_bready[4]),
.m4_arid(rtl_m_arid[4]), .m4_araddr(rtl_m_araddr[4]), .m4_arlen(rtl_m_arlen[4]),
.m4_arsize(rtl_m_arsize[4]), .m4_arburst(rtl_m_arburst[4]), .m4_arlock(rtl_m_arlock[4]),
.m4_arcache(rtl_m_arcache[4]), .m4_arprot(rtl_m_arprot[4]), .m4_arqos(rtl_m_arqos[4]),
.m4_arvalid(rtl_m_arvalid[4]), .m4_arready(rtl_m_arready[4]),
.m4_rid(rtl_m_rid[4]), .m4_rdata(rtl_m_rdata[4]), .m4_rresp(rtl_m_rresp[4]),
.m4_rlast(rtl_m_rlast[4]), .m4_rvalid(rtl_m_rvalid[4]), .m4_rready(rtl_m_rready[4]),

// Master 5 connections
.m5_awid(rtl_m_awid[5]), .m5_awaddr(rtl_m_awaddr[5]), .m5_awlen(rtl_m_awlen[5]),
.m5_awsize(rtl_m_awsize[5]), .m5_awburst(rtl_m_awburst[5]), .m5_awlock(rtl_m_awlock[5]),
.m5_awcache(rtl_m_awcache[5]), .m5_awprot(rtl_m_awprot[5]), .m5_awqos(rtl_m_awqos[5]),
.m5_awvalid(rtl_m_awvalid[5]), .m5_awready(rtl_m_awready[5]),
.m5_wdata(rtl_m_wdata[5]), .m5_wstrb(rtl_m_wstrb[5]), .m5_wlast(rtl_m_wlast[5]),
.m5_wvalid(rtl_m_wvalid[5]), .m5_wready(rtl_m_wready[5]),
.m5_bid(rtl_m_bid[5]), .m5_bresp(rtl_m_bresp[5]), .m5_bvalid(rtl_m_bvalid[5]), .m5_bready(rtl_m_bready[5]),
.m5_arid(rtl_m_arid[5]), .m5_araddr(rtl_m_araddr[5]), .m5_arlen(rtl_m_arlen[5]),
.m5_arsize(rtl_m_arsize[5]), .m5_arburst(rtl_m_arburst[5]), .m5_arlock(rtl_m_arlock[5]),
.m5_arcache(rtl_m_arcache[5]), .m5_arprot(rtl_m_arprot[5]), .m5_arqos(rtl_m_arqos[5]),
.m5_arvalid(rtl_m_arvalid[5]), .m5_arready(rtl_m_arready[5]),
.m5_rid(rtl_m_rid[5]), .m5_rdata(rtl_m_rdata[5]), .m5_rresp(rtl_m_rresp[5]),
.m5_rlast(rtl_m_rlast[5]), .m5_rvalid(rtl_m_rvalid[5]), .m5_rready(rtl_m_rready[5]),

// Master 6 connections
.m6_awid(rtl_m_awid[6]), .m6_awaddr(rtl_m_awaddr[6]), .m6_awlen(rtl_m_awlen[6]),
.m6_awsize(rtl_m_awsize[6]), .m6_awburst(rtl_m_awburst[6]), .m6_awlock(rtl_m_awlock[6]),
.m6_awcache(rtl_m_awcache[6]), .m6_awprot(rtl_m_awprot[6]), .m6_awqos(rtl_m_awqos[6]),
.m6_awvalid(rtl_m_awvalid[6]), .m6_awready(rtl_m_awready[6]),
.m6_wdata(rtl_m_wdata[6]), .m6_wstrb(rtl_m_wstrb[6]), .m6_wlast(rtl_m_wlast[6]),
.m6_wvalid(rtl_m_wvalid[6]), .m6_wready(rtl_m_wready[6]),
.m6_bid(rtl_m_bid[6]), .m6_bresp(rtl_m_bresp[6]), .m6_bvalid(rtl_m_bvalid[6]), .m6_bready(rtl_m_bready[6]),
.m6_arid(rtl_m_arid[6]), .m6_araddr(rtl_m_araddr[6]), .m6_arlen(rtl_m_arlen[6]),
.m6_arsize(rtl_m_arsize[6]), .m6_arburst(rtl_m_arburst[6]), .m6_arlock(rtl_m_arlock[6]),
.m6_arcache(rtl_m_arcache[6]), .m6_arprot(rtl_m_arprot[6]), .m6_arqos(rtl_m_arqos[6]),
.m6_arvalid(rtl_m_arvalid[6]), .m6_arready(rtl_m_arready[6]),
.m6_rid(rtl_m_rid[6]), .m6_rdata(rtl_m_rdata[6]), .m6_rresp(rtl_m_rresp[6]),
.m6_rlast(rtl_m_rlast[6]), .m6_rvalid(rtl_m_rvalid[6]), .m6_rready(rtl_m_rready[6]),

// Master 7 connections
.m7_awid(rtl_m_awid[7]), .m7_awaddr(rtl_m_awaddr[7]), .m7_awlen(rtl_m_awlen[7]),
.m7_awsize(rtl_m_awsize[7]), .m7_awburst(rtl_m_awburst[7]), .m7_awlock(rtl_m_awlock[7]),
.m7_awcache(rtl_m_awcache[7]), .m7_awprot(rtl_m_awprot[7]), .m7_awqos(rtl_m_awqos[7]),
.m7_awvalid(rtl_m_awvalid[7]), .m7_awready(rtl_m_awready[7]),
.m7_wdata(rtl_m_wdata[7]), .m7_wstrb(rtl_m_wstrb[7]), .m7_wlast(rtl_m_wlast[7]),
.m7_wvalid(rtl_m_wvalid[7]), .m7_wready(rtl_m_wready[7]),
.m7_bid(rtl_m_bid[7]), .m7_bresp(rtl_m_bresp[7]), .m7_bvalid(rtl_m_bvalid[7]), .m7_bready(rtl_m_bready[7]),
.m7_arid(rtl_m_arid[7]), .m7_araddr(rtl_m_araddr[7]), .m7_arlen(rtl_m_arlen[7]),
.m7_arsize(rtl_m_arsize[7]), .m7_arburst(rtl_m_arburst[7]), .m7_arlock(rtl_m_arlock[7]),
.m7_arcache(rtl_m_arcache[7]), .m7_arprot(rtl_m_arprot[7]), .m7_arqos(rtl_m_arqos[7]),
.m7_arvalid(rtl_m_arvalid[7]), .m7_arready(rtl_m_arready[7]),
.m7_rid(rtl_m_rid[7]), .m7_rdata(rtl_m_rdata[7]), .m7_rresp(rtl_m_rresp[7]),
.m7_rlast(rtl_m_rlast[7]), .m7_rvalid(rtl_m_rvalid[7]), .m7_rready(rtl_m_rready[7]),

// Master 8 connections
.m8_awid(rtl_m_awid[8]), .m8_awaddr(rtl_m_awaddr[8]), .m8_awlen(rtl_m_awlen[8]),
.m8_awsize(rtl_m_awsize[8]), .m8_awburst(rtl_m_awburst[8]), .m8_awlock(rtl_m_awlock[8]),
.m8_awcache(rtl_m_awcache[8]), .m8_awprot(rtl_m_awprot[8]), .m8_awqos(rtl_m_awqos[8]),
.m8_awvalid(rtl_m_awvalid[8]), .m8_awready(rtl_m_awready[8]),
.m8_wdata(rtl_m_wdata[8]), .m8_wstrb(rtl_m_wstrb[8]), .m8_wlast(rtl_m_wlast[8]),
.m8_wvalid(rtl_m_wvalid[8]), .m8_wready(rtl_m_wready[8]),
.m8_bid(rtl_m_bid[8]), .m8_bresp(rtl_m_bresp[8]), .m8_bvalid(rtl_m_bvalid[8]), .m8_bready(rtl_m_bready[8]),
.m8_arid(rtl_m_arid[8]), .m8_araddr(rtl_m_araddr[8]), .m8_arlen(rtl_m_arlen[8]),
.m8_arsize(rtl_m_arsize[8]), .m8_arburst(rtl_m_arburst[8]), .m8_arlock(rtl_m_arlock[8]),
.m8_arcache(rtl_m_arcache[8]), .m8_arprot(rtl_m_arprot[8]), .m8_arqos(rtl_m_arqos[8]),
.m8_arvalid(rtl_m_arvalid[8]), .m8_arready(rtl_m_arready[8]),
.m8_rid(rtl_m_rid[8]), .m8_rdata(rtl_m_rdata[8]), .m8_rresp(rtl_m_rresp[8]),
.m8_rlast(rtl_m_rlast[8]), .m8_rvalid(rtl_m_rvalid[8]), .m8_rready(rtl_m_rready[8]),

// Master 9 connections
.m9_awid(rtl_m_awid[9]), .m9_awaddr(rtl_m_awaddr[9]), .m9_awlen(rtl_m_awlen[9]),
.m9_awsize(rtl_m_awsize[9]), .m9_awburst(rtl_m_awburst[9]), .m9_awlock(rtl_m_awlock[9]),
.m9_awcache(rtl_m_awcache[9]), .m9_awprot(rtl_m_awprot[9]), .m9_awqos(rtl_m_awqos[9]),
.m9_awvalid(rtl_m_awvalid[9]), .m9_awready(rtl_m_awready[9]),
.m9_wdata(rtl_m_wdata[9]), .m9_wstrb(rtl_m_wstrb[9]), .m9_wlast(rtl_m_wlast[9]),
.m9_wvalid(rtl_m_wvalid[9]), .m9_wready(rtl_m_wready[9]),
.m9_bid(rtl_m_bid[9]), .m9_bresp(rtl_m_bresp[9]), .m9_bvalid(rtl_m_bvalid[9]), .m9_bready(rtl_m_bready[9]),
.m9_arid(rtl_m_arid[9]), .m9_araddr(rtl_m_araddr[9]), .m9_arlen(rtl_m_arlen[9]),
.m9_arsize(rtl_m_arsize[9]), .m9_arburst(rtl_m_arburst[9]), .m9_arlock(rtl_m_arlock[9]),
.m9_arcache(rtl_m_arcache[9]), .m9_arprot(rtl_m_arprot[9]), .m9_arqos(rtl_m_arqos[9]),
.m9_arvalid(rtl_m_arvalid[9]), .m9_arready(rtl_m_arready[9]),
.m9_rid(rtl_m_rid[9]), .m9_rdata(rtl_m_rdata[9]), .m9_rresp(rtl_m_rresp[9]),
.m9_rlast(rtl_m_rlast[9]), .m9_rvalid(rtl_m_rvalid[9]), .m9_rready(rtl_m_rready[9]),

// Master 10 connections
.m10_awid(rtl_m_awid[10]), .m10_awaddr(rtl_m_awaddr[10]), .m10_awlen(rtl_m_awlen[10]),
.m10_awsize(rtl_m_awsize[10]), .m10_awburst(rtl_m_awburst[10]), .m10_awlock(rtl_m_awlock[10]),
.m10_awcache(rtl_m_awcache[10]), .m10_awprot(rtl_m_awprot[10]), .m10_awqos(rtl_m_awqos[10]),
.m10_awvalid(rtl_m_awvalid[10]), .m10_awready(rtl_m_awready[10]),
.m10_wdata(rtl_m_wdata[10]), .m10_wstrb(rtl_m_wstrb[10]), .m10_wlast(rtl_m_wlast[10]),
.m10_wvalid(rtl_m_wvalid[10]), .m10_wready(rtl_m_wready[10]),
.m10_bid(rtl_m_bid[10]), .m10_bresp(rtl_m_bresp[10]), .m10_bvalid(rtl_m_bvalid[10]), .m10_bready(rtl_m_bready[10]),
.m10_arid(rtl_m_arid[10]), .m10_araddr(rtl_m_araddr[10]), .m10_arlen(rtl_m_arlen[10]),
.m10_arsize(rtl_m_arsize[10]), .m10_arburst(rtl_m_arburst[10]), .m10_arlock(rtl_m_arlock[10]),
.m10_arcache(rtl_m_arcache[10]), .m10_arprot(rtl_m_arprot[10]), .m10_arqos(rtl_m_arqos[10]),
.m10_arvalid(rtl_m_arvalid[10]), .m10_arready(rtl_m_arready[10]),
.m10_rid(rtl_m_rid[10]), .m10_rdata(rtl_m_rdata[10]), .m10_rresp(rtl_m_rresp[10]),
.m10_rlast(rtl_m_rlast[10]), .m10_rvalid(rtl_m_rvalid[10]), .m10_rready(rtl_m_rready[10]),

// Master 11 connections
.m11_awid(rtl_m_awid[11]), .m11_awaddr(rtl_m_awaddr[11]), .m11_awlen(rtl_m_awlen[11]),
.m11_awsize(rtl_m_awsize[11]), .m11_awburst(rtl_m_awburst[11]), .m11_awlock(rtl_m_awlock[11]),
.m11_awcache(rtl_m_awcache[11]), .m11_awprot(rtl_m_awprot[11]), .m11_awqos(rtl_m_awqos[11]),
.m11_awvalid(rtl_m_awvalid[11]), .m11_awready(rtl_m_awready[11]),
.m11_wdata(rtl_m_wdata[11]), .m11_wstrb(rtl_m_wstrb[11]), .m11_wlast(rtl_m_wlast[11]),
.m11_wvalid(rtl_m_wvalid[11]), .m11_wready(rtl_m_wready[11]),
.m11_bid(rtl_m_bid[11]), .m11_bresp(rtl_m_bresp[11]), .m11_bvalid(rtl_m_bvalid[11]), .m11_bready(rtl_m_bready[11]),
.m11_arid(rtl_m_arid[11]), .m11_araddr(rtl_m_araddr[11]), .m11_arlen(rtl_m_arlen[11]),
.m11_arsize(rtl_m_arsize[11]), .m11_arburst(rtl_m_arburst[11]), .m11_arlock(rtl_m_arlock[11]),
.m11_arcache(rtl_m_arcache[11]), .m11_arprot(rtl_m_arprot[11]), .m11_arqos(rtl_m_arqos[11]),
.m11_arvalid(rtl_m_arvalid[11]), .m11_arready(rtl_m_arready[11]),
.m11_rid(rtl_m_rid[11]), .m11_rdata(rtl_m_rdata[11]), .m11_rresp(rtl_m_rresp[11]),
.m11_rlast(rtl_m_rlast[11]), .m11_rvalid(rtl_m_rvalid[11]), .m11_rready(rtl_m_rready[11]),

// Master 12 connections
.m12_awid(rtl_m_awid[12]), .m12_awaddr(rtl_m_awaddr[12]), .m12_awlen(rtl_m_awlen[12]),
.m12_awsize(rtl_m_awsize[12]), .m12_awburst(rtl_m_awburst[12]), .m12_awlock(rtl_m_awlock[12]),
.m12_awcache(rtl_m_awcache[12]), .m12_awprot(rtl_m_awprot[12]), .m12_awqos(rtl_m_awqos[12]),
.m12_awvalid(rtl_m_awvalid[12]), .m12_awready(rtl_m_awready[12]),
.m12_wdata(rtl_m_wdata[12]), .m12_wstrb(rtl_m_wstrb[12]), .m12_wlast(rtl_m_wlast[12]),
.m12_wvalid(rtl_m_wvalid[12]), .m12_wready(rtl_m_wready[12]),
.m12_bid(rtl_m_bid[12]), .m12_bresp(rtl_m_bresp[12]), .m12_bvalid(rtl_m_bvalid[12]), .m12_bready(rtl_m_bready[12]),
.m12_arid(rtl_m_arid[12]), .m12_araddr(rtl_m_araddr[12]), .m12_arlen(rtl_m_arlen[12]),
.m12_arsize(rtl_m_arsize[12]), .m12_arburst(rtl_m_arburst[12]), .m12_arlock(rtl_m_arlock[12]),
.m12_arcache(rtl_m_arcache[12]), .m12_arprot(rtl_m_arprot[12]), .m12_arqos(rtl_m_arqos[12]),
.m12_arvalid(rtl_m_arvalid[12]), .m12_arready(rtl_m_arready[12]),
.m12_rid(rtl_m_rid[12]), .m12_rdata(rtl_m_rdata[12]), .m12_rresp(rtl_m_rresp[12]),
.m12_rlast(rtl_m_rlast[12]), .m12_rvalid(rtl_m_rvalid[12]), .m12_rready(rtl_m_rready[12]),

// Master 13 connections
.m13_awid(rtl_m_awid[13]), .m13_awaddr(rtl_m_awaddr[13]), .m13_awlen(rtl_m_awlen[13]),
.m13_awsize(rtl_m_awsize[13]), .m13_awburst(rtl_m_awburst[13]), .m13_awlock(rtl_m_awlock[13]),
.m13_awcache(rtl_m_awcache[13]), .m13_awprot(rtl_m_awprot[13]), .m13_awqos(rtl_m_awqos[13]),
.m13_awvalid(rtl_m_awvalid[13]), .m13_awready(rtl_m_awready[13]),
.m13_wdata(rtl_m_wdata[13]), .m13_wstrb(rtl_m_wstrb[13]), .m13_wlast(rtl_m_wlast[13]),
.m13_wvalid(rtl_m_wvalid[13]), .m13_wready(rtl_m_wready[13]),
.m13_bid(rtl_m_bid[13]), .m13_bresp(rtl_m_bresp[13]), .m13_bvalid(rtl_m_bvalid[13]), .m13_bready(rtl_m_bready[13]),
.m13_arid(rtl_m_arid[13]), .m13_araddr(rtl_m_araddr[13]), .m13_arlen(rtl_m_arlen[13]),
.m13_arsize(rtl_m_arsize[13]), .m13_arburst(rtl_m_arburst[13]), .m13_arlock(rtl_m_arlock[13]),
.m13_arcache(rtl_m_arcache[13]), .m13_arprot(rtl_m_arprot[13]), .m13_arqos(rtl_m_arqos[13]),
.m13_arvalid(rtl_m_arvalid[13]), .m13_arready(rtl_m_arready[13]),
.m13_rid(rtl_m_rid[13]), .m13_rdata(rtl_m_rdata[13]), .m13_rresp(rtl_m_rresp[13]),
.m13_rlast(rtl_m_rlast[13]), .m13_rvalid(rtl_m_rvalid[13]), .m13_rready(rtl_m_rready[13]),

// Master 14 connections
.m14_awid(rtl_m_awid[14]), .m14_awaddr(rtl_m_awaddr[14]), .m14_awlen(rtl_m_awlen[14]),
.m14_awsize(rtl_m_awsize[14]), .m14_awburst(rtl_m_awburst[14]), .m14_awlock(rtl_m_awlock[14]),
.m14_awcache(rtl_m_awcache[14]), .m14_awprot(rtl_m_awprot[14]), .m14_awqos(rtl_m_awqos[14]),
.m14_awvalid(rtl_m_awvalid[14]), .m14_awready(rtl_m_awready[14]),
.m14_wdata(rtl_m_wdata[14]), .m14_wstrb(rtl_m_wstrb[14]), .m14_wlast(rtl_m_wlast[14]),
.m14_wvalid(rtl_m_wvalid[14]), .m14_wready(rtl_m_wready[14]),
.m14_bid(rtl_m_bid[14]), .m14_bresp(rtl_m_bresp[14]), .m14_bvalid(rtl_m_bvalid[14]), .m14_bready(rtl_m_bready[14]),
.m14_arid(rtl_m_arid[14]), .m14_araddr(rtl_m_araddr[14]), .m14_arlen(rtl_m_arlen[14]),
.m14_arsize(rtl_m_arsize[14]), .m14_arburst(rtl_m_arburst[14]), .m14_arlock(rtl_m_arlock[14]),
.m14_arcache(rtl_m_arcache[14]), .m14_arprot(rtl_m_arprot[14]), .m14_arqos(rtl_m_arqos[14]),
.m14_arvalid(rtl_m_arvalid[14]), .m14_arready(rtl_m_arready[14]),
.m14_rid(rtl_m_rid[14]), .m14_rdata(rtl_m_rdata[14]), .m14_rresp(rtl_m_rresp[14]),
.m14_rlast(rtl_m_rlast[14]), .m14_rvalid(rtl_m_rvalid[14]), .m14_rready(rtl_m_rready[14]),

// Slave 1 connections
.s1_awid(rtl_s_awid[1]), .s1_awaddr(rtl_s_awaddr[1]), .s1_awlen(rtl_s_awlen[1]),
.s1_awsize(rtl_s_awsize[1]), .s1_awburst(rtl_s_awburst[1]), .s1_awlock(rtl_s_awlock[1]),
.s1_awcache(rtl_s_awcache[1]), .s1_awprot(rtl_s_awprot[1]), .s1_awqos(rtl_s_awqos[1]),
.s1_awvalid(rtl_s_awvalid[1]), .s1_awready(rtl_s_awready[1]),
.s1_wdata(rtl_s_wdata[1]), .s1_wstrb(rtl_s_wstrb[1]), .s1_wlast(rtl_s_wlast[1]),
.s1_wvalid(rtl_s_wvalid[1]), .s1_wready(rtl_s_wready[1]),
.s1_bid(rtl_s_bid[1]), .s1_bresp(rtl_s_bresp[1]), .s1_bvalid(rtl_s_bvalid[1]), .s1_bready(rtl_s_bready[1]),
.s1_arid(rtl_s_arid[1]), .s1_araddr(rtl_s_araddr[1]), .s1_arlen(rtl_s_arlen[1]),
.s1_arsize(rtl_s_arsize[1]), .s1_arburst(rtl_s_arburst[1]), .s1_arlock(rtl_s_arlock[1]),
.s1_arcache(rtl_s_arcache[1]), .s1_arprot(rtl_s_arprot[1]), .s1_arqos(rtl_s_arqos[1]),
.s1_arvalid(rtl_s_arvalid[1]), .s1_arready(rtl_s_arready[1]),
.s1_rid(rtl_s_rid[1]), .s1_rdata(rtl_s_rdata[1]), .s1_rresp(rtl_s_rresp[1]),
.s1_rlast(rtl_s_rlast[1]), .s1_rvalid(rtl_s_rvalid[1]), .s1_rready(rtl_s_rready[1]),

// Slave 2 connections
.s2_awid(rtl_s_awid[2]), .s2_awaddr(rtl_s_awaddr[2]), .s2_awlen(rtl_s_awlen[2]),
.s2_awsize(rtl_s_awsize[2]), .s2_awburst(rtl_s_awburst[2]), .s2_awlock(rtl_s_awlock[2]),
.s2_awcache(rtl_s_awcache[2]), .s2_awprot(rtl_s_awprot[2]), .s2_awqos(rtl_s_awqos[2]),
.s2_awvalid(rtl_s_awvalid[2]), .s2_awready(rtl_s_awready[2]),
.s2_wdata(rtl_s_wdata[2]), .s2_wstrb(rtl_s_wstrb[2]), .s2_wlast(rtl_s_wlast[2]),
.s2_wvalid(rtl_s_wvalid[2]), .s2_wready(rtl_s_wready[2]),
.s2_bid(rtl_s_bid[2]), .s2_bresp(rtl_s_bresp[2]), .s2_bvalid(rtl_s_bvalid[2]), .s2_bready(rtl_s_bready[2]),
.s2_arid(rtl_s_arid[2]), .s2_araddr(rtl_s_araddr[2]), .s2_arlen(rtl_s_arlen[2]),
.s2_arsize(rtl_s_arsize[2]), .s2_arburst(rtl_s_arburst[2]), .s2_arlock(rtl_s_arlock[2]),
.s2_arcache(rtl_s_arcache[2]), .s2_arprot(rtl_s_arprot[2]), .s2_arqos(rtl_s_arqos[2]),
.s2_arvalid(rtl_s_arvalid[2]), .s2_arready(rtl_s_arready[2]),
.s2_rid(rtl_s_rid[2]), .s2_rdata(rtl_s_rdata[2]), .s2_rresp(rtl_s_rresp[2]),
.s2_rlast(rtl_s_rlast[2]), .s2_rvalid(rtl_s_rvalid[2]), .s2_rready(rtl_s_rready[2]),

// Slave 3 connections
.s3_awid(rtl_s_awid[3]), .s3_awaddr(rtl_s_awaddr[3]), .s3_awlen(rtl_s_awlen[3]),
.s3_awsize(rtl_s_awsize[3]), .s3_awburst(rtl_s_awburst[3]), .s3_awlock(rtl_s_awlock[3]),
.s3_awcache(rtl_s_awcache[3]), .s3_awprot(rtl_s_awprot[3]), .s3_awqos(rtl_s_awqos[3]),
.s3_awvalid(rtl_s_awvalid[3]), .s3_awready(rtl_s_awready[3]),
.s3_wdata(rtl_s_wdata[3]), .s3_wstrb(rtl_s_wstrb[3]), .s3_wlast(rtl_s_wlast[3]),
.s3_wvalid(rtl_s_wvalid[3]), .s3_wready(rtl_s_wready[3]),
.s3_bid(rtl_s_bid[3]), .s3_bresp(rtl_s_bresp[3]), .s3_bvalid(rtl_s_bvalid[3]), .s3_bready(rtl_s_bready[3]),
.s3_arid(rtl_s_arid[3]), .s3_araddr(rtl_s_araddr[3]), .s3_arlen(rtl_s_arlen[3]),
.s3_arsize(rtl_s_arsize[3]), .s3_arburst(rtl_s_arburst[3]), .s3_arlock(rtl_s_arlock[3]),
.s3_arcache(rtl_s_arcache[3]), .s3_arprot(rtl_s_arprot[3]), .s3_arqos(rtl_s_arqos[3]),
.s3_arvalid(rtl_s_arvalid[3]), .s3_arready(rtl_s_arready[3]),
.s3_rid(rtl_s_rid[3]), .s3_rdata(rtl_s_rdata[3]), .s3_rresp(rtl_s_rresp[3]),
.s3_rlast(rtl_s_rlast[3]), .s3_rvalid(rtl_s_rvalid[3]), .s3_rready(rtl_s_rready[3]),

// Slave 4 connections
.s4_awid(rtl_s_awid[4]), .s4_awaddr(rtl_s_awaddr[4]), .s4_awlen(rtl_s_awlen[4]),
.s4_awsize(rtl_s_awsize[4]), .s4_awburst(rtl_s_awburst[4]), .s4_awlock(rtl_s_awlock[4]),
.s4_awcache(rtl_s_awcache[4]), .s4_awprot(rtl_s_awprot[4]), .s4_awqos(rtl_s_awqos[4]),
.s4_awvalid(rtl_s_awvalid[4]), .s4_awready(rtl_s_awready[4]),
.s4_wdata(rtl_s_wdata[4]), .s4_wstrb(rtl_s_wstrb[4]), .s4_wlast(rtl_s_wlast[4]),
.s4_wvalid(rtl_s_wvalid[4]), .s4_wready(rtl_s_wready[4]),
.s4_bid(rtl_s_bid[4]), .s4_bresp(rtl_s_bresp[4]), .s4_bvalid(rtl_s_bvalid[4]), .s4_bready(rtl_s_bready[4]),
.s4_arid(rtl_s_arid[4]), .s4_araddr(rtl_s_araddr[4]), .s4_arlen(rtl_s_arlen[4]),
.s4_arsize(rtl_s_arsize[4]), .s4_arburst(rtl_s_arburst[4]), .s4_arlock(rtl_s_arlock[4]),
.s4_arcache(rtl_s_arcache[4]), .s4_arprot(rtl_s_arprot[4]), .s4_arqos(rtl_s_arqos[4]),
.s4_arvalid(rtl_s_arvalid[4]), .s4_arready(rtl_s_arready[4]),
.s4_rid(rtl_s_rid[4]), .s4_rdata(rtl_s_rdata[4]), .s4_rresp(rtl_s_rresp[4]),
.s4_rlast(rtl_s_rlast[4]), .s4_rvalid(rtl_s_rvalid[4]), .s4_rready(rtl_s_rready[4]),

// Slave 5 connections
.s5_awid(rtl_s_awid[5]), .s5_awaddr(rtl_s_awaddr[5]), .s5_awlen(rtl_s_awlen[5]),
.s5_awsize(rtl_s_awsize[5]), .s5_awburst(rtl_s_awburst[5]), .s5_awlock(rtl_s_awlock[5]),
.s5_awcache(rtl_s_awcache[5]), .s5_awprot(rtl_s_awprot[5]), .s5_awqos(rtl_s_awqos[5]),
.s5_awvalid(rtl_s_awvalid[5]), .s5_awready(rtl_s_awready[5]),
.s5_wdata(rtl_s_wdata[5]), .s5_wstrb(rtl_s_wstrb[5]), .s5_wlast(rtl_s_wlast[5]),
.s5_wvalid(rtl_s_wvalid[5]), .s5_wready(rtl_s_wready[5]),
.s5_bid(rtl_s_bid[5]), .s5_bresp(rtl_s_bresp[5]), .s5_bvalid(rtl_s_bvalid[5]), .s5_bready(rtl_s_bready[5]),
.s5_arid(rtl_s_arid[5]), .s5_araddr(rtl_s_araddr[5]), .s5_arlen(rtl_s_arlen[5]),
.s5_arsize(rtl_s_arsize[5]), .s5_arburst(rtl_s_arburst[5]), .s5_arlock(rtl_s_arlock[5]),
.s5_arcache(rtl_s_arcache[5]), .s5_arprot(rtl_s_arprot[5]), .s5_arqos(rtl_s_arqos[5]),
.s5_arvalid(rtl_s_arvalid[5]), .s5_arready(rtl_s_arready[5]),
.s5_rid(rtl_s_rid[5]), .s5_rdata(rtl_s_rdata[5]), .s5_rresp(rtl_s_rresp[5]),
.s5_rlast(rtl_s_rlast[5]), .s5_rvalid(rtl_s_rvalid[5]), .s5_rready(rtl_s_rready[5]),

// Slave 6 connections
.s6_awid(rtl_s_awid[6]), .s6_awaddr(rtl_s_awaddr[6]), .s6_awlen(rtl_s_awlen[6]),
.s6_awsize(rtl_s_awsize[6]), .s6_awburst(rtl_s_awburst[6]), .s6_awlock(rtl_s_awlock[6]),
.s6_awcache(rtl_s_awcache[6]), .s6_awprot(rtl_s_awprot[6]), .s6_awqos(rtl_s_awqos[6]),
.s6_awvalid(rtl_s_awvalid[6]), .s6_awready(rtl_s_awready[6]),
.s6_wdata(rtl_s_wdata[6]), .s6_wstrb(rtl_s_wstrb[6]), .s6_wlast(rtl_s_wlast[6]),
.s6_wvalid(rtl_s_wvalid[6]), .s6_wready(rtl_s_wready[6]),
.s6_bid(rtl_s_bid[6]), .s6_bresp(rtl_s_bresp[6]), .s6_bvalid(rtl_s_bvalid[6]), .s6_bready(rtl_s_bready[6]),
.s6_arid(rtl_s_arid[6]), .s6_araddr(rtl_s_araddr[6]), .s6_arlen(rtl_s_arlen[6]),
.s6_arsize(rtl_s_arsize[6]), .s6_arburst(rtl_s_arburst[6]), .s6_arlock(rtl_s_arlock[6]),
.s6_arcache(rtl_s_arcache[6]), .s6_arprot(rtl_s_arprot[6]), .s6_arqos(rtl_s_arqos[6]),
.s6_arvalid(rtl_s_arvalid[6]), .s6_arready(rtl_s_arready[6]),
.s6_rid(rtl_s_rid[6]), .s6_rdata(rtl_s_rdata[6]), .s6_rresp(rtl_s_rresp[6]),
.s6_rlast(rtl_s_rlast[6]), .s6_rvalid(rtl_s_rvalid[6]), .s6_rready(rtl_s_rready[6]),

// Slave 7 connections
.s7_awid(rtl_s_awid[7]), .s7_awaddr(rtl_s_awaddr[7]), .s7_awlen(rtl_s_awlen[7]),
.s7_awsize(rtl_s_awsize[7]), .s7_awburst(rtl_s_awburst[7]), .s7_awlock(rtl_s_awlock[7]),
.s7_awcache(rtl_s_awcache[7]), .s7_awprot(rtl_s_awprot[7]), .s7_awqos(rtl_s_awqos[7]),
.s7_awvalid(rtl_s_awvalid[7]), .s7_awready(rtl_s_awready[7]),
.s7_wdata(rtl_s_wdata[7]), .s7_wstrb(rtl_s_wstrb[7]), .s7_wlast(rtl_s_wlast[7]),
.s7_wvalid(rtl_s_wvalid[7]), .s7_wready(rtl_s_wready[7]),
.s7_bid(rtl_s_bid[7]), .s7_bresp(rtl_s_bresp[7]), .s7_bvalid(rtl_s_bvalid[7]), .s7_bready(rtl_s_bready[7]),
.s7_arid(rtl_s_arid[7]), .s7_araddr(rtl_s_araddr[7]), .s7_arlen(rtl_s_arlen[7]),
.s7_arsize(rtl_s_arsize[7]), .s7_arburst(rtl_s_arburst[7]), .s7_arlock(rtl_s_arlock[7]),
.s7_arcache(rtl_s_arcache[7]), .s7_arprot(rtl_s_arprot[7]), .s7_arqos(rtl_s_arqos[7]),
.s7_arvalid(rtl_s_arvalid[7]), .s7_arready(rtl_s_arready[7]),
.s7_rid(rtl_s_rid[7]), .s7_rdata(rtl_s_rdata[7]), .s7_rresp(rtl_s_rresp[7]),
.s7_rlast(rtl_s_rlast[7]), .s7_rvalid(rtl_s_rvalid[7]), .s7_rready(rtl_s_rready[7]),

// Slave 8 connections
.s8_awid(rtl_s_awid[8]), .s8_awaddr(rtl_s_awaddr[8]), .s8_awlen(rtl_s_awlen[8]),
.s8_awsize(rtl_s_awsize[8]), .s8_awburst(rtl_s_awburst[8]), .s8_awlock(rtl_s_awlock[8]),
.s8_awcache(rtl_s_awcache[8]), .s8_awprot(rtl_s_awprot[8]), .s8_awqos(rtl_s_awqos[8]),
.s8_awvalid(rtl_s_awvalid[8]), .s8_awready(rtl_s_awready[8]),
.s8_wdata(rtl_s_wdata[8]), .s8_wstrb(rtl_s_wstrb[8]), .s8_wlast(rtl_s_wlast[8]),
.s8_wvalid(rtl_s_wvalid[8]), .s8_wready(rtl_s_wready[8]),
.s8_bid(rtl_s_bid[8]), .s8_bresp(rtl_s_bresp[8]), .s8_bvalid(rtl_s_bvalid[8]), .s8_bready(rtl_s_bready[8]),
.s8_arid(rtl_s_arid[8]), .s8_araddr(rtl_s_araddr[8]), .s8_arlen(rtl_s_arlen[8]),
.s8_arsize(rtl_s_arsize[8]), .s8_arburst(rtl_s_arburst[8]), .s8_arlock(rtl_s_arlock[8]),
.s8_arcache(rtl_s_arcache[8]), .s8_arprot(rtl_s_arprot[8]), .s8_arqos(rtl_s_arqos[8]),
.s8_arvalid(rtl_s_arvalid[8]), .s8_arready(rtl_s_arready[8]),
.s8_rid(rtl_s_rid[8]), .s8_rdata(rtl_s_rdata[8]), .s8_rresp(rtl_s_rresp[8]),
.s8_rlast(rtl_s_rlast[8]), .s8_rvalid(rtl_s_rvalid[8]), .s8_rready(rtl_s_rready[8]),

// Slave 9 connections
.s9_awid(rtl_s_awid[9]), .s9_awaddr(rtl_s_awaddr[9]), .s9_awlen(rtl_s_awlen[9]),
.s9_awsize(rtl_s_awsize[9]), .s9_awburst(rtl_s_awburst[9]), .s9_awlock(rtl_s_awlock[9]),
.s9_awcache(rtl_s_awcache[9]), .s9_awprot(rtl_s_awprot[9]), .s9_awqos(rtl_s_awqos[9]),
.s9_awvalid(rtl_s_awvalid[9]), .s9_awready(rtl_s_awready[9]),
.s9_wdata(rtl_s_wdata[9]), .s9_wstrb(rtl_s_wstrb[9]), .s9_wlast(rtl_s_wlast[9]),
.s9_wvalid(rtl_s_wvalid[9]), .s9_wready(rtl_s_wready[9]),
.s9_bid(rtl_s_bid[9]), .s9_bresp(rtl_s_bresp[9]), .s9_bvalid(rtl_s_bvalid[9]), .s9_bready(rtl_s_bready[9]),
.s9_arid(rtl_s_arid[9]), .s9_araddr(rtl_s_araddr[9]), .s9_arlen(rtl_s_arlen[9]),
.s9_arsize(rtl_s_arsize[9]), .s9_arburst(rtl_s_arburst[9]), .s9_arlock(rtl_s_arlock[9]),
.s9_arcache(rtl_s_arcache[9]), .s9_arprot(rtl_s_arprot[9]), .s9_arqos(rtl_s_arqos[9]),
.s9_arvalid(rtl_s_arvalid[9]), .s9_arready(rtl_s_arready[9]),
.s9_rid(rtl_s_rid[9]), .s9_rdata(rtl_s_rdata[9]), .s9_rresp(rtl_s_rresp[9]),
.s9_rlast(rtl_s_rlast[9]), .s9_rvalid(rtl_s_rvalid[9]), .s9_rready(rtl_s_rready[9]),

// Slave 10 connections
.s10_awid(rtl_s_awid[10]), .s10_awaddr(rtl_s_awaddr[10]), .s10_awlen(rtl_s_awlen[10]),
.s10_awsize(rtl_s_awsize[10]), .s10_awburst(rtl_s_awburst[10]), .s10_awlock(rtl_s_awlock[10]),
.s10_awcache(rtl_s_awcache[10]), .s10_awprot(rtl_s_awprot[10]), .s10_awqos(rtl_s_awqos[10]),
.s10_awvalid(rtl_s_awvalid[10]), .s10_awready(rtl_s_awready[10]),
.s10_wdata(rtl_s_wdata[10]), .s10_wstrb(rtl_s_wstrb[10]), .s10_wlast(rtl_s_wlast[10]),
.s10_wvalid(rtl_s_wvalid[10]), .s10_wready(rtl_s_wready[10]),
.s10_bid(rtl_s_bid[10]), .s10_bresp(rtl_s_bresp[10]), .s10_bvalid(rtl_s_bvalid[10]), .s10_bready(rtl_s_bready[10]),
.s10_arid(rtl_s_arid[10]), .s10_araddr(rtl_s_araddr[10]), .s10_arlen(rtl_s_arlen[10]),
.s10_arsize(rtl_s_arsize[10]), .s10_arburst(rtl_s_arburst[10]), .s10_arlock(rtl_s_arlock[10]),
.s10_arcache(rtl_s_arcache[10]), .s10_arprot(rtl_s_arprot[10]), .s10_arqos(rtl_s_arqos[10]),
.s10_arvalid(rtl_s_arvalid[10]), .s10_arready(rtl_s_arready[10]),
.s10_rid(rtl_s_rid[10]), .s10_rdata(rtl_s_rdata[10]), .s10_rresp(rtl_s_rresp[10]),
.s10_rlast(rtl_s_rlast[10]), .s10_rvalid(rtl_s_rvalid[10]), .s10_rready(rtl_s_rready[10]),

// Slave 11 connections
.s11_awid(rtl_s_awid[11]), .s11_awaddr(rtl_s_awaddr[11]), .s11_awlen(rtl_s_awlen[11]),
.s11_awsize(rtl_s_awsize[11]), .s11_awburst(rtl_s_awburst[11]), .s11_awlock(rtl_s_awlock[11]),
.s11_awcache(rtl_s_awcache[11]), .s11_awprot(rtl_s_awprot[11]), .s11_awqos(rtl_s_awqos[11]),
.s11_awvalid(rtl_s_awvalid[11]), .s11_awready(rtl_s_awready[11]),
.s11_wdata(rtl_s_wdata[11]), .s11_wstrb(rtl_s_wstrb[11]), .s11_wlast(rtl_s_wlast[11]),
.s11_wvalid(rtl_s_wvalid[11]), .s11_wready(rtl_s_wready[11]),
.s11_bid(rtl_s_bid[11]), .s11_bresp(rtl_s_bresp[11]), .s11_bvalid(rtl_s_bvalid[11]), .s11_bready(rtl_s_bready[11]),
.s11_arid(rtl_s_arid[11]), .s11_araddr(rtl_s_araddr[11]), .s11_arlen(rtl_s_arlen[11]),
.s11_arsize(rtl_s_arsize[11]), .s11_arburst(rtl_s_arburst[11]), .s11_arlock(rtl_s_arlock[11]),
.s11_arcache(rtl_s_arcache[11]), .s11_arprot(rtl_s_arprot[11]), .s11_arqos(rtl_s_arqos[11]),
.s11_arvalid(rtl_s_arvalid[11]), .s11_arready(rtl_s_arready[11]),
.s11_rid(rtl_s_rid[11]), .s11_rdata(rtl_s_rdata[11]), .s11_rresp(rtl_s_rresp[11]),
.s11_rlast(rtl_s_rlast[11]), .s11_rvalid(rtl_s_rvalid[11]), .s11_rready(rtl_s_rready[11]),

// Slave 12 connections
.s12_awid(rtl_s_awid[12]), .s12_awaddr(rtl_s_awaddr[12]), .s12_awlen(rtl_s_awlen[12]),
.s12_awsize(rtl_s_awsize[12]), .s12_awburst(rtl_s_awburst[12]), .s12_awlock(rtl_s_awlock[12]),
.s12_awcache(rtl_s_awcache[12]), .s12_awprot(rtl_s_awprot[12]), .s12_awqos(rtl_s_awqos[12]),
.s12_awvalid(rtl_s_awvalid[12]), .s12_awready(rtl_s_awready[12]),
.s12_wdata(rtl_s_wdata[12]), .s12_wstrb(rtl_s_wstrb[12]), .s12_wlast(rtl_s_wlast[12]),
.s12_wvalid(rtl_s_wvalid[12]), .s12_wready(rtl_s_wready[12]),
.s12_bid(rtl_s_bid[12]), .s12_bresp(rtl_s_bresp[12]), .s12_bvalid(rtl_s_bvalid[12]), .s12_bready(rtl_s_bready[12]),
.s12_arid(rtl_s_arid[12]), .s12_araddr(rtl_s_araddr[12]), .s12_arlen(rtl_s_arlen[12]),
.s12_arsize(rtl_s_arsize[12]), .s12_arburst(rtl_s_arburst[12]), .s12_arlock(rtl_s_arlock[12]),
.s12_arcache(rtl_s_arcache[12]), .s12_arprot(rtl_s_arprot[12]), .s12_arqos(rtl_s_arqos[12]),
.s12_arvalid(rtl_s_arvalid[12]), .s12_arready(rtl_s_arready[12]),
.s12_rid(rtl_s_rid[12]), .s12_rdata(rtl_s_rdata[12]), .s12_rresp(rtl_s_rresp[12]),
.s12_rlast(rtl_s_rlast[12]), .s12_rvalid(rtl_s_rvalid[12]), .s12_rready(rtl_s_rready[12]),

// Slave 13 connections
.s13_awid(rtl_s_awid[13]), .s13_awaddr(rtl_s_awaddr[13]), .s13_awlen(rtl_s_awlen[13]),
.s13_awsize(rtl_s_awsize[13]), .s13_awburst(rtl_s_awburst[13]), .s13_awlock(rtl_s_awlock[13]),
.s13_awcache(rtl_s_awcache[13]), .s13_awprot(rtl_s_awprot[13]), .s13_awqos(rtl_s_awqos[13]),
.s13_awvalid(rtl_s_awvalid[13]), .s13_awready(rtl_s_awready[13]),
.s13_wdata(rtl_s_wdata[13]), .s13_wstrb(rtl_s_wstrb[13]), .s13_wlast(rtl_s_wlast[13]),
.s13_wvalid(rtl_s_wvalid[13]), .s13_wready(rtl_s_wready[13]),
.s13_bid(rtl_s_bid[13]), .s13_bresp(rtl_s_bresp[13]), .s13_bvalid(rtl_s_bvalid[13]), .s13_bready(rtl_s_bready[13]),
.s13_arid(rtl_s_arid[13]), .s13_araddr(rtl_s_araddr[13]), .s13_arlen(rtl_s_arlen[13]),
.s13_arsize(rtl_s_arsize[13]), .s13_arburst(rtl_s_arburst[13]), .s13_arlock(rtl_s_arlock[13]),
.s13_arcache(rtl_s_arcache[13]), .s13_arprot(rtl_s_arprot[13]), .s13_arqos(rtl_s_arqos[13]),
.s13_arvalid(rtl_s_arvalid[13]), .s13_arready(rtl_s_arready[13]),
.s13_rid(rtl_s_rid[13]), .s13_rdata(rtl_s_rdata[13]), .s13_rresp(rtl_s_rresp[13]),
.s13_rlast(rtl_s_rlast[13]), .s13_rvalid(rtl_s_rvalid[13]), .s13_rready(rtl_s_rready[13]),

// Slave 14 connections
.s14_awid(rtl_s_awid[14]), .s14_awaddr(rtl_s_awaddr[14]), .s14_awlen(rtl_s_awlen[14]),
.s14_awsize(rtl_s_awsize[14]), .s14_awburst(rtl_s_awburst[14]), .s14_awlock(rtl_s_awlock[14]),
.s14_awcache(rtl_s_awcache[14]), .s14_awprot(rtl_s_awprot[14]), .s14_awqos(rtl_s_awqos[14]),
.s14_awvalid(rtl_s_awvalid[14]), .s14_awready(rtl_s_awready[14]),
.s14_wdata(rtl_s_wdata[14]), .s14_wstrb(rtl_s_wstrb[14]), .s14_wlast(rtl_s_wlast[14]),
.s14_wvalid(rtl_s_wvalid[14]), .s14_wready(rtl_s_wready[14]),
.s14_bid(rtl_s_bid[14]), .s14_bresp(rtl_s_bresp[14]), .s14_bvalid(rtl_s_bvalid[14]), .s14_bready(rtl_s_bready[14]),
.s14_arid(rtl_s_arid[14]), .s14_araddr(rtl_s_araddr[14]), .s14_arlen(rtl_s_arlen[14]),
.s14_arsize(rtl_s_arsize[14]), .s14_arburst(rtl_s_arburst[14]), .s14_arlock(rtl_s_arlock[14]),
.s14_arcache(rtl_s_arcache[14]), .s14_arprot(rtl_s_arprot[14]), .s14_arqos(rtl_s_arqos[14]),
.s14_arvalid(rtl_s_arvalid[14]), .s14_arready(rtl_s_arready[14]),
.s14_rid(rtl_s_rid[14]), .s14_rdata(rtl_s_rdata[14]), .s14_rresp(rtl_s_rresp[14]),
.s14_rlast(rtl_s_rlast[14]), .s14_rvalid(rtl_s_rvalid[14]), .s14_rready(rtl_s_rready[14])