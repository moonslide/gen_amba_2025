// Stub slave monitor BFM - replace with actual implementation  
interface axi4_slave_monitor_bfm(input aclk, input aresetn);
endinterface
