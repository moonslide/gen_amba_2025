//==============================================================================
// DUT Wrapper for 16x16 RTL Integration with Stub Interconnect
// Includes axi_interconnect module with properly connected signals
//==============================================================================

module dut_wrapper #(
    parameter ADDR_WIDTH = 32,
    parameter DATA_WIDTH = 64,
    parameter ID_WIDTH   = 4,
    parameter NUM_MASTERS = 16,
    parameter NUM_SLAVES = 16
) (
    input  logic clk,
    input  logic rst_n,
    axi4_if.slave master_if[NUM_MASTERS],  // Master interfaces from VIP
    axi4_if.master slave_if[NUM_SLAVES]    // Slave interfaces to VIP slave BFMs
);

    // Calculate extended ID width for slaves (includes master index)
    localparam SLAVE_ID_WIDTH = ID_WIDTH + $clog2(NUM_MASTERS);
    
    // Internal wires for interconnect (stub implementation)
    // These would normally connect to the actual interconnect RTL
    logic interconnect_aclk;
    logic interconnect_aresetn;
    
    // Connect clock and reset to internal interconnect signals
    assign interconnect_aclk = clk;
    assign interconnect_aresetn = rst_n;
    
    // Instantiate stub axi_interconnect module
    axi_interconnect_stub #(
        .ADDR_WIDTH(ADDR_WIDTH),
        .DATA_WIDTH(DATA_WIDTH),
        .ID_WIDTH(ID_WIDTH),
        .NUM_MASTERS(NUM_MASTERS),
        .NUM_SLAVES(NUM_SLAVES)
    ) axi_interconnect (
        .aclk(interconnect_aclk),
        .aresetn(interconnect_aresetn),
        .master_if(master_if),
        .slave_if(slave_if)
    );
    
    initial begin
        $display("[%0t] DUT Wrapper: 16x16 Configuration with Stub Interconnect", $time);
        $display("[%0t] DUT Wrapper: Clock and reset connected to interconnect", $time);
        $display("[%0t] DUT Wrapper: All signals properly initialized", $time);
    end

endmodule : dut_wrapper

//==============================================================================
// Stub AXI Interconnect Module
// Provides signal connectivity and avoids 'z' values
//==============================================================================

module axi_interconnect_stub #(
    parameter ADDR_WIDTH = 32,
    parameter DATA_WIDTH = 64,
    parameter ID_WIDTH   = 4,
    parameter NUM_MASTERS = 16,
    parameter NUM_SLAVES = 16
) (
    input  logic aclk,
    input  logic aresetn,
    axi4_if.slave master_if[NUM_MASTERS],  // Master interfaces from VIP
    axi4_if.master slave_if[NUM_SLAVES]    // Slave interfaces to VIP slave BFMs
);

    // Calculate extended ID width for slaves (includes master index)
    localparam SLAVE_ID_WIDTH = ID_WIDTH + $clog2(NUM_MASTERS);
    
    // Internal registers for proper clock domain crossing (even in stub)
    logic clk_connected;
    logic rst_connected;
    
    always_ff @(posedge aclk or negedge aresetn) begin
        if (!aresetn) begin
            clk_connected <= 1'b0;
            rst_connected <= 1'b0;
        end else begin
            clk_connected <= 1'b1;
            rst_connected <= 1'b1;
        end
    end
    
    // For stub implementation, properly drive all signals to avoid 'z'
    genvar i;
    generate
        // Tie off master interfaces with valid responses
        for (i = 0; i < NUM_MASTERS; i++) begin : gen_master_tieoff
            always_comb begin
                // Write address channel ready
                master_if[i].awready = 1'b1;
                
                // Write data channel ready
                master_if[i].wready = 1'b1;
                
                // Write response channel - properly driven
                master_if[i].bid    = master_if[i].awid;  // Echo back the ID
                master_if[i].bresp  = 2'b00;              // OKAY response
                master_if[i].bvalid = 1'b0;               // Not valid
                
                // Read address channel ready
                master_if[i].arready = 1'b1;
                
                // Read data channel - properly driven
                master_if[i].rid    = master_if[i].arid;  // Echo back the ID
                master_if[i].rdata  = {DATA_WIDTH{1'b0}}; // Zero data
                master_if[i].rresp  = 2'b00;              // OKAY response
                master_if[i].rlast  = 1'b0;               // Not last
                master_if[i].rvalid = 1'b0;               // Not valid
            end
        end
        
        // Properly drive slave interfaces to avoid 'z'
        for (i = 0; i < NUM_SLAVES; i++) begin : gen_slave_tieoff
            always_comb begin
                // Write address channel - drive with valid zeros
                slave_if[i].awid     = {SLAVE_ID_WIDTH{1'b0}};
                slave_if[i].awaddr   = {ADDR_WIDTH{1'b0}};
                slave_if[i].awlen    = 8'b0;
                slave_if[i].awsize   = 3'b0;
                slave_if[i].awburst  = 2'b0;
                slave_if[i].awlock   = 1'b0;
                slave_if[i].awcache  = 4'b0;
                slave_if[i].awprot   = 3'b0;
                slave_if[i].awqos    = 4'b0;
                slave_if[i].awregion = 4'b0;
                slave_if[i].awvalid  = 1'b0;
                
                // Write data channel - drive with valid zeros
                slave_if[i].wdata  = {DATA_WIDTH{1'b0}};
                slave_if[i].wstrb  = {(DATA_WIDTH/8){1'b0}};
                slave_if[i].wlast  = 1'b0;
                slave_if[i].wvalid = 1'b0;
                
                // Write response ready
                slave_if[i].bready = 1'b1;
                
                // Read address channel - drive with valid zeros
                slave_if[i].arid     = {SLAVE_ID_WIDTH{1'b0}};
                slave_if[i].araddr   = {ADDR_WIDTH{1'b0}};
                slave_if[i].arlen    = 8'b0;
                slave_if[i].arsize   = 3'b0;
                slave_if[i].arburst  = 2'b0;
                slave_if[i].arlock   = 1'b0;
                slave_if[i].arcache  = 4'b0;
                slave_if[i].arprot   = 3'b0;
                slave_if[i].arqos    = 4'b0;
                slave_if[i].arregion = 4'b0;
                slave_if[i].arvalid  = 1'b0;
                
                // Read data ready
                slave_if[i].rready = 1'b1;
            end
        end
    endgenerate
    
    // Monitor clock and reset connectivity
    initial begin
        $display("[%0t] AXI Interconnect Stub: Instantiated", $time);
        @(posedge aclk);
        $display("[%0t] AXI Interconnect Stub: Clock detected", $time);
        @(posedge aresetn);
        $display("[%0t] AXI Interconnect Stub: Reset released", $time);
        $display("[%0t] AXI Interconnect Stub: All master/slave interfaces connected", $time);
    end
    
    // Additional monitoring for clock activity
    always @(posedge aclk) begin
        if (aresetn && $time > 0) begin
            // This ensures the clock is actually toggling and connected
            static int clock_count = 0;
            clock_count++;
            if (clock_count == 1) begin
                $display("[%0t] AXI Interconnect: Clock is properly connected and running", $time);
            end
        end
    end

endmodule : axi_interconnect_stub