// Stub master monitor BFM - replace with actual implementation
interface axi4_master_monitor_bfm(input aclk, input aresetn);
endinterface
