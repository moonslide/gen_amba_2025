// Slave wire declarations for Slaves 1-14
// This file is included in dut_wrapper_real_rtl.sv
// Note: RTL outputs ID_WIDTH=4, but slaves need SLAVE_ID_WIDTH (includes master index)

// Slave 1
wire [RTL_ID_WIDTH-1:0]     s1_awid;
wire [ADDR_WIDTH-1:0]       s1_awaddr;
wire [7:0]                  s1_awlen;
wire [2:0]                  s1_awsize;
wire [1:0]                  s1_awburst;
wire                        s1_awlock;
wire [3:0]                  s1_awcache;
wire [2:0]                  s1_awprot;
wire [3:0]                  s1_awqos;
wire                        s1_awvalid;
wire                        s1_awready;
wire [DATA_WIDTH-1:0]       s1_wdata;
wire [DATA_WIDTH/8-1:0]     s1_wstrb;
wire                        s1_wlast;
wire                        s1_wvalid;
wire                        s1_wready;
wire [RTL_ID_WIDTH-1:0]     s1_bid;
wire [1:0]                  s1_bresp;
wire                        s1_bvalid;
wire                        s1_bready;
wire [RTL_ID_WIDTH-1:0]     s1_arid;
wire [ADDR_WIDTH-1:0]       s1_araddr;
wire [7:0]                  s1_arlen;
wire [2:0]                  s1_arsize;
wire [1:0]                  s1_arburst;
wire                        s1_arlock;
wire [3:0]                  s1_arcache;
wire [2:0]                  s1_arprot;
wire [3:0]                  s1_arqos;
wire                        s1_arvalid;
wire                        s1_arready;
wire [RTL_ID_WIDTH-1:0]     s1_rid;
wire [DATA_WIDTH-1:0]       s1_rdata;
wire [1:0]                  s1_rresp;
wire                        s1_rlast;
wire                        s1_rvalid;
wire                        s1_rready;

// Slave 2
wire [RTL_ID_WIDTH-1:0]     s2_awid;
wire [ADDR_WIDTH-1:0]       s2_awaddr;
wire [7:0]                  s2_awlen;
wire [2:0]                  s2_awsize;
wire [1:0]                  s2_awburst;
wire                        s2_awlock;
wire [3:0]                  s2_awcache;
wire [2:0]                  s2_awprot;
wire [3:0]                  s2_awqos;
wire                        s2_awvalid;
wire                        s2_awready;
wire [DATA_WIDTH-1:0]       s2_wdata;
wire [DATA_WIDTH/8-1:0]     s2_wstrb;
wire                        s2_wlast;
wire                        s2_wvalid;
wire                        s2_wready;
wire [RTL_ID_WIDTH-1:0]     s2_bid;
wire [1:0]                  s2_bresp;
wire                        s2_bvalid;
wire                        s2_bready;
wire [RTL_ID_WIDTH-1:0]     s2_arid;
wire [ADDR_WIDTH-1:0]       s2_araddr;
wire [7:0]                  s2_arlen;
wire [2:0]                  s2_arsize;
wire [1:0]                  s2_arburst;
wire                        s2_arlock;
wire [3:0]                  s2_arcache;
wire [2:0]                  s2_arprot;
wire [3:0]                  s2_arqos;
wire                        s2_arvalid;
wire                        s2_arready;
wire [RTL_ID_WIDTH-1:0]     s2_rid;
wire [DATA_WIDTH-1:0]       s2_rdata;
wire [1:0]                  s2_rresp;
wire                        s2_rlast;
wire                        s2_rvalid;
wire                        s2_rready;

// Slave 3
wire [RTL_ID_WIDTH-1:0]     s3_awid;
wire [ADDR_WIDTH-1:0]       s3_awaddr;
wire [7:0]                  s3_awlen;
wire [2:0]                  s3_awsize;
wire [1:0]                  s3_awburst;
wire                        s3_awlock;
wire [3:0]                  s3_awcache;
wire [2:0]                  s3_awprot;
wire [3:0]                  s3_awqos;
wire                        s3_awvalid;
wire                        s3_awready;
wire [DATA_WIDTH-1:0]       s3_wdata;
wire [DATA_WIDTH/8-1:0]     s3_wstrb;
wire                        s3_wlast;
wire                        s3_wvalid;
wire                        s3_wready;
wire [RTL_ID_WIDTH-1:0]     s3_bid;
wire [1:0]                  s3_bresp;
wire                        s3_bvalid;
wire                        s3_bready;
wire [RTL_ID_WIDTH-1:0]     s3_arid;
wire [ADDR_WIDTH-1:0]       s3_araddr;
wire [7:0]                  s3_arlen;
wire [2:0]                  s3_arsize;
wire [1:0]                  s3_arburst;
wire                        s3_arlock;
wire [3:0]                  s3_arcache;
wire [2:0]                  s3_arprot;
wire [3:0]                  s3_arqos;
wire                        s3_arvalid;
wire                        s3_arready;
wire [RTL_ID_WIDTH-1:0]     s3_rid;
wire [DATA_WIDTH-1:0]       s3_rdata;
wire [1:0]                  s3_rresp;
wire                        s3_rlast;
wire                        s3_rvalid;
wire                        s3_rready;

// Slave 4
wire [RTL_ID_WIDTH-1:0]     s4_awid;
wire [ADDR_WIDTH-1:0]       s4_awaddr;
wire [7:0]                  s4_awlen;
wire [2:0]                  s4_awsize;
wire [1:0]                  s4_awburst;
wire                        s4_awlock;
wire [3:0]                  s4_awcache;
wire [2:0]                  s4_awprot;
wire [3:0]                  s4_awqos;
wire                        s4_awvalid;
wire                        s4_awready;
wire [DATA_WIDTH-1:0]       s4_wdata;
wire [DATA_WIDTH/8-1:0]     s4_wstrb;
wire                        s4_wlast;
wire                        s4_wvalid;
wire                        s4_wready;
wire [RTL_ID_WIDTH-1:0]     s4_bid;
wire [1:0]                  s4_bresp;
wire                        s4_bvalid;
wire                        s4_bready;
wire [RTL_ID_WIDTH-1:0]     s4_arid;
wire [ADDR_WIDTH-1:0]       s4_araddr;
wire [7:0]                  s4_arlen;
wire [2:0]                  s4_arsize;
wire [1:0]                  s4_arburst;
wire                        s4_arlock;
wire [3:0]                  s4_arcache;
wire [2:0]                  s4_arprot;
wire [3:0]                  s4_arqos;
wire                        s4_arvalid;
wire                        s4_arready;
wire [RTL_ID_WIDTH-1:0]     s4_rid;
wire [DATA_WIDTH-1:0]       s4_rdata;
wire [1:0]                  s4_rresp;
wire                        s4_rlast;
wire                        s4_rvalid;
wire                        s4_rready;

// Slave 5
wire [RTL_ID_WIDTH-1:0]     s5_awid;
wire [ADDR_WIDTH-1:0]       s5_awaddr;
wire [7:0]                  s5_awlen;
wire [2:0]                  s5_awsize;
wire [1:0]                  s5_awburst;
wire                        s5_awlock;
wire [3:0]                  s5_awcache;
wire [2:0]                  s5_awprot;
wire [3:0]                  s5_awqos;
wire                        s5_awvalid;
wire                        s5_awready;
wire [DATA_WIDTH-1:0]       s5_wdata;
wire [DATA_WIDTH/8-1:0]     s5_wstrb;
wire                        s5_wlast;
wire                        s5_wvalid;
wire                        s5_wready;
wire [RTL_ID_WIDTH-1:0]     s5_bid;
wire [1:0]                  s5_bresp;
wire                        s5_bvalid;
wire                        s5_bready;
wire [RTL_ID_WIDTH-1:0]     s5_arid;
wire [ADDR_WIDTH-1:0]       s5_araddr;
wire [7:0]                  s5_arlen;
wire [2:0]                  s5_arsize;
wire [1:0]                  s5_arburst;
wire                        s5_arlock;
wire [3:0]                  s5_arcache;
wire [2:0]                  s5_arprot;
wire [3:0]                  s5_arqos;
wire                        s5_arvalid;
wire                        s5_arready;
wire [RTL_ID_WIDTH-1:0]     s5_rid;
wire [DATA_WIDTH-1:0]       s5_rdata;
wire [1:0]                  s5_rresp;
wire                        s5_rlast;
wire                        s5_rvalid;
wire                        s5_rready;

// Slave 6
wire [RTL_ID_WIDTH-1:0]     s6_awid;
wire [ADDR_WIDTH-1:0]       s6_awaddr;
wire [7:0]                  s6_awlen;
wire [2:0]                  s6_awsize;
wire [1:0]                  s6_awburst;
wire                        s6_awlock;
wire [3:0]                  s6_awcache;
wire [2:0]                  s6_awprot;
wire [3:0]                  s6_awqos;
wire                        s6_awvalid;
wire                        s6_awready;
wire [DATA_WIDTH-1:0]       s6_wdata;
wire [DATA_WIDTH/8-1:0]     s6_wstrb;
wire                        s6_wlast;
wire                        s6_wvalid;
wire                        s6_wready;
wire [RTL_ID_WIDTH-1:0]     s6_bid;
wire [1:0]                  s6_bresp;
wire                        s6_bvalid;
wire                        s6_bready;
wire [RTL_ID_WIDTH-1:0]     s6_arid;
wire [ADDR_WIDTH-1:0]       s6_araddr;
wire [7:0]                  s6_arlen;
wire [2:0]                  s6_arsize;
wire [1:0]                  s6_arburst;
wire                        s6_arlock;
wire [3:0]                  s6_arcache;
wire [2:0]                  s6_arprot;
wire [3:0]                  s6_arqos;
wire                        s6_arvalid;
wire                        s6_arready;
wire [RTL_ID_WIDTH-1:0]     s6_rid;
wire [DATA_WIDTH-1:0]       s6_rdata;
wire [1:0]                  s6_rresp;
wire                        s6_rlast;
wire                        s6_rvalid;
wire                        s6_rready;

// Slave 7
wire [RTL_ID_WIDTH-1:0]     s7_awid;
wire [ADDR_WIDTH-1:0]       s7_awaddr;
wire [7:0]                  s7_awlen;
wire [2:0]                  s7_awsize;
wire [1:0]                  s7_awburst;
wire                        s7_awlock;
wire [3:0]                  s7_awcache;
wire [2:0]                  s7_awprot;
wire [3:0]                  s7_awqos;
wire                        s7_awvalid;
wire                        s7_awready;
wire [DATA_WIDTH-1:0]       s7_wdata;
wire [DATA_WIDTH/8-1:0]     s7_wstrb;
wire                        s7_wlast;
wire                        s7_wvalid;
wire                        s7_wready;
wire [RTL_ID_WIDTH-1:0]     s7_bid;
wire [1:0]                  s7_bresp;
wire                        s7_bvalid;
wire                        s7_bready;
wire [RTL_ID_WIDTH-1:0]     s7_arid;
wire [ADDR_WIDTH-1:0]       s7_araddr;
wire [7:0]                  s7_arlen;
wire [2:0]                  s7_arsize;
wire [1:0]                  s7_arburst;
wire                        s7_arlock;
wire [3:0]                  s7_arcache;
wire [2:0]                  s7_arprot;
wire [3:0]                  s7_arqos;
wire                        s7_arvalid;
wire                        s7_arready;
wire [RTL_ID_WIDTH-1:0]     s7_rid;
wire [DATA_WIDTH-1:0]       s7_rdata;
wire [1:0]                  s7_rresp;
wire                        s7_rlast;
wire                        s7_rvalid;
wire                        s7_rready;

// Slave 8
wire [RTL_ID_WIDTH-1:0]     s8_awid;
wire [ADDR_WIDTH-1:0]       s8_awaddr;
wire [7:0]                  s8_awlen;
wire [2:0]                  s8_awsize;
wire [1:0]                  s8_awburst;
wire                        s8_awlock;
wire [3:0]                  s8_awcache;
wire [2:0]                  s8_awprot;
wire [3:0]                  s8_awqos;
wire                        s8_awvalid;
wire                        s8_awready;
wire [DATA_WIDTH-1:0]       s8_wdata;
wire [DATA_WIDTH/8-1:0]     s8_wstrb;
wire                        s8_wlast;
wire                        s8_wvalid;
wire                        s8_wready;
wire [RTL_ID_WIDTH-1:0]     s8_bid;
wire [1:0]                  s8_bresp;
wire                        s8_bvalid;
wire                        s8_bready;
wire [RTL_ID_WIDTH-1:0]     s8_arid;
wire [ADDR_WIDTH-1:0]       s8_araddr;
wire [7:0]                  s8_arlen;
wire [2:0]                  s8_arsize;
wire [1:0]                  s8_arburst;
wire                        s8_arlock;
wire [3:0]                  s8_arcache;
wire [2:0]                  s8_arprot;
wire [3:0]                  s8_arqos;
wire                        s8_arvalid;
wire                        s8_arready;
wire [RTL_ID_WIDTH-1:0]     s8_rid;
wire [DATA_WIDTH-1:0]       s8_rdata;
wire [1:0]                  s8_rresp;
wire                        s8_rlast;
wire                        s8_rvalid;
wire                        s8_rready;

// Slave 9
wire [RTL_ID_WIDTH-1:0]     s9_awid;
wire [ADDR_WIDTH-1:0]       s9_awaddr;
wire [7:0]                  s9_awlen;
wire [2:0]                  s9_awsize;
wire [1:0]                  s9_awburst;
wire                        s9_awlock;
wire [3:0]                  s9_awcache;
wire [2:0]                  s9_awprot;
wire [3:0]                  s9_awqos;
wire                        s9_awvalid;
wire                        s9_awready;
wire [DATA_WIDTH-1:0]       s9_wdata;
wire [DATA_WIDTH/8-1:0]     s9_wstrb;
wire                        s9_wlast;
wire                        s9_wvalid;
wire                        s9_wready;
wire [RTL_ID_WIDTH-1:0]     s9_bid;
wire [1:0]                  s9_bresp;
wire                        s9_bvalid;
wire                        s9_bready;
wire [RTL_ID_WIDTH-1:0]     s9_arid;
wire [ADDR_WIDTH-1:0]       s9_araddr;
wire [7:0]                  s9_arlen;
wire [2:0]                  s9_arsize;
wire [1:0]                  s9_arburst;
wire                        s9_arlock;
wire [3:0]                  s9_arcache;
wire [2:0]                  s9_arprot;
wire [3:0]                  s9_arqos;
wire                        s9_arvalid;
wire                        s9_arready;
wire [RTL_ID_WIDTH-1:0]     s9_rid;
wire [DATA_WIDTH-1:0]       s9_rdata;
wire [1:0]                  s9_rresp;
wire                        s9_rlast;
wire                        s9_rvalid;
wire                        s9_rready;

// Slave 10
wire [RTL_ID_WIDTH-1:0]     s10_awid;
wire [ADDR_WIDTH-1:0]       s10_awaddr;
wire [7:0]                  s10_awlen;
wire [2:0]                  s10_awsize;
wire [1:0]                  s10_awburst;
wire                        s10_awlock;
wire [3:0]                  s10_awcache;
wire [2:0]                  s10_awprot;
wire [3:0]                  s10_awqos;
wire                        s10_awvalid;
wire                        s10_awready;
wire [DATA_WIDTH-1:0]       s10_wdata;
wire [DATA_WIDTH/8-1:0]     s10_wstrb;
wire                        s10_wlast;
wire                        s10_wvalid;
wire                        s10_wready;
wire [RTL_ID_WIDTH-1:0]     s10_bid;
wire [1:0]                  s10_bresp;
wire                        s10_bvalid;
wire                        s10_bready;
wire [RTL_ID_WIDTH-1:0]     s10_arid;
wire [ADDR_WIDTH-1:0]       s10_araddr;
wire [7:0]                  s10_arlen;
wire [2:0]                  s10_arsize;
wire [1:0]                  s10_arburst;
wire                        s10_arlock;
wire [3:0]                  s10_arcache;
wire [2:0]                  s10_arprot;
wire [3:0]                  s10_arqos;
wire                        s10_arvalid;
wire                        s10_arready;
wire [RTL_ID_WIDTH-1:0]     s10_rid;
wire [DATA_WIDTH-1:0]       s10_rdata;
wire [1:0]                  s10_rresp;
wire                        s10_rlast;
wire                        s10_rvalid;
wire                        s10_rready;

// Slave 11
wire [RTL_ID_WIDTH-1:0]     s11_awid;
wire [ADDR_WIDTH-1:0]       s11_awaddr;
wire [7:0]                  s11_awlen;
wire [2:0]                  s11_awsize;
wire [1:0]                  s11_awburst;
wire                        s11_awlock;
wire [3:0]                  s11_awcache;
wire [2:0]                  s11_awprot;
wire [3:0]                  s11_awqos;
wire                        s11_awvalid;
wire                        s11_awready;
wire [DATA_WIDTH-1:0]       s11_wdata;
wire [DATA_WIDTH/8-1:0]     s11_wstrb;
wire                        s11_wlast;
wire                        s11_wvalid;
wire                        s11_wready;
wire [RTL_ID_WIDTH-1:0]     s11_bid;
wire [1:0]                  s11_bresp;
wire                        s11_bvalid;
wire                        s11_bready;
wire [RTL_ID_WIDTH-1:0]     s11_arid;
wire [ADDR_WIDTH-1:0]       s11_araddr;
wire [7:0]                  s11_arlen;
wire [2:0]                  s11_arsize;
wire [1:0]                  s11_arburst;
wire                        s11_arlock;
wire [3:0]                  s11_arcache;
wire [2:0]                  s11_arprot;
wire [3:0]                  s11_arqos;
wire                        s11_arvalid;
wire                        s11_arready;
wire [RTL_ID_WIDTH-1:0]     s11_rid;
wire [DATA_WIDTH-1:0]       s11_rdata;
wire [1:0]                  s11_rresp;
wire                        s11_rlast;
wire                        s11_rvalid;
wire                        s11_rready;

// Slave 12
wire [RTL_ID_WIDTH-1:0]     s12_awid;
wire [ADDR_WIDTH-1:0]       s12_awaddr;
wire [7:0]                  s12_awlen;
wire [2:0]                  s12_awsize;
wire [1:0]                  s12_awburst;
wire                        s12_awlock;
wire [3:0]                  s12_awcache;
wire [2:0]                  s12_awprot;
wire [3:0]                  s12_awqos;
wire                        s12_awvalid;
wire                        s12_awready;
wire [DATA_WIDTH-1:0]       s12_wdata;
wire [DATA_WIDTH/8-1:0]     s12_wstrb;
wire                        s12_wlast;
wire                        s12_wvalid;
wire                        s12_wready;
wire [RTL_ID_WIDTH-1:0]     s12_bid;
wire [1:0]                  s12_bresp;
wire                        s12_bvalid;
wire                        s12_bready;
wire [RTL_ID_WIDTH-1:0]     s12_arid;
wire [ADDR_WIDTH-1:0]       s12_araddr;
wire [7:0]                  s12_arlen;
wire [2:0]                  s12_arsize;
wire [1:0]                  s12_arburst;
wire                        s12_arlock;
wire [3:0]                  s12_arcache;
wire [2:0]                  s12_arprot;
wire [3:0]                  s12_arqos;
wire                        s12_arvalid;
wire                        s12_arready;
wire [RTL_ID_WIDTH-1:0]     s12_rid;
wire [DATA_WIDTH-1:0]       s12_rdata;
wire [1:0]                  s12_rresp;
wire                        s12_rlast;
wire                        s12_rvalid;
wire                        s12_rready;

// Slave 13
wire [RTL_ID_WIDTH-1:0]     s13_awid;
wire [ADDR_WIDTH-1:0]       s13_awaddr;
wire [7:0]                  s13_awlen;
wire [2:0]                  s13_awsize;
wire [1:0]                  s13_awburst;
wire                        s13_awlock;
wire [3:0]                  s13_awcache;
wire [2:0]                  s13_awprot;
wire [3:0]                  s13_awqos;
wire                        s13_awvalid;
wire                        s13_awready;
wire [DATA_WIDTH-1:0]       s13_wdata;
wire [DATA_WIDTH/8-1:0]     s13_wstrb;
wire                        s13_wlast;
wire                        s13_wvalid;
wire                        s13_wready;
wire [RTL_ID_WIDTH-1:0]     s13_bid;
wire [1:0]                  s13_bresp;
wire                        s13_bvalid;
wire                        s13_bready;
wire [RTL_ID_WIDTH-1:0]     s13_arid;
wire [ADDR_WIDTH-1:0]       s13_araddr;
wire [7:0]                  s13_arlen;
wire [2:0]                  s13_arsize;
wire [1:0]                  s13_arburst;
wire                        s13_arlock;
wire [3:0]                  s13_arcache;
wire [2:0]                  s13_arprot;
wire [3:0]                  s13_arqos;
wire                        s13_arvalid;
wire                        s13_arready;
wire [RTL_ID_WIDTH-1:0]     s13_rid;
wire [DATA_WIDTH-1:0]       s13_rdata;
wire [1:0]                  s13_rresp;
wire                        s13_rlast;
wire                        s13_rvalid;
wire                        s13_rready;

// Slave 14
wire [RTL_ID_WIDTH-1:0]     s14_awid;
wire [ADDR_WIDTH-1:0]       s14_awaddr;
wire [7:0]                  s14_awlen;
wire [2:0]                  s14_awsize;
wire [1:0]                  s14_awburst;
wire                        s14_awlock;
wire [3:0]                  s14_awcache;
wire [2:0]                  s14_awprot;
wire [3:0]                  s14_awqos;
wire                        s14_awvalid;
wire                        s14_awready;
wire [DATA_WIDTH-1:0]       s14_wdata;
wire [DATA_WIDTH/8-1:0]     s14_wstrb;
wire                        s14_wlast;
wire                        s14_wvalid;
wire                        s14_wready;
wire [RTL_ID_WIDTH-1:0]     s14_bid;
wire [1:0]                  s14_bresp;
wire                        s14_bvalid;
wire                        s14_bready;
wire [RTL_ID_WIDTH-1:0]     s14_arid;
wire [ADDR_WIDTH-1:0]       s14_araddr;
wire [7:0]                  s14_arlen;
wire [2:0]                  s14_arsize;
wire [1:0]                  s14_arburst;
wire                        s14_arlock;
wire [3:0]                  s14_arcache;
wire [2:0]                  s14_arprot;
wire [3:0]                  s14_arqos;
wire                        s14_arvalid;
wire                        s14_arready;
wire [RTL_ID_WIDTH-1:0]     s14_rid;
wire [DATA_WIDTH-1:0]       s14_rdata;
wire [1:0]                  s14_rresp;
wire                        s14_rlast;
wire                        s14_rvalid;
wire                        s14_rready;