        // Master 1 connections
        .m1_awid(m1_awid),
        .m1_awaddr(m1_awaddr),
        .m1_awlen(m1_awlen),
        .m1_awsize(m1_awsize),
        .m1_awburst(m1_awburst),
        .m1_awlock(m1_awlock),
        .m1_awcache(m1_awcache),
        .m1_awprot(m1_awprot),
        .m1_awqos(m1_awqos),
        .m1_awvalid(m1_awvalid),
        .m1_awready(m1_awready),
        .m1_wdata(m1_wdata),
        .m1_wstrb(m1_wstrb),
        .m1_wlast(m1_wlast),
        .m1_wvalid(m1_wvalid),
        .m1_wready(m1_wready),
        .m1_bid(m1_bid),
        .m1_bresp(m1_bresp),
        .m1_bvalid(m1_bvalid),
        .m1_bready(m1_bready),
        .m1_arid(m1_arid),
        .m1_araddr(m1_araddr),
        .m1_arlen(m1_arlen),
        .m1_arsize(m1_arsize),
        .m1_arburst(m1_arburst),
        .m1_arlock(m1_arlock),
        .m1_arcache(m1_arcache),
        .m1_arprot(m1_arprot),
        .m1_arqos(m1_arqos),
        .m1_arvalid(m1_arvalid),
        .m1_arready(m1_arready),
        .m1_rid(m1_rid),
        .m1_rdata(m1_rdata),
        .m1_rresp(m1_rresp),
        .m1_rlast(m1_rlast),
        .m1_rvalid(m1_rvalid),
        .m1_rready(m1_rready),
        // Master 2 connections
        .m2_awid(m2_awid),
        .m2_awaddr(m2_awaddr),
        .m2_awlen(m2_awlen),
        .m2_awsize(m2_awsize),
        .m2_awburst(m2_awburst),
        .m2_awlock(m2_awlock),
        .m2_awcache(m2_awcache),
        .m2_awprot(m2_awprot),
        .m2_awqos(m2_awqos),
        .m2_awvalid(m2_awvalid),
        .m2_awready(m2_awready),
        .m2_wdata(m2_wdata),
        .m2_wstrb(m2_wstrb),
        .m2_wlast(m2_wlast),
        .m2_wvalid(m2_wvalid),
        .m2_wready(m2_wready),
        .m2_bid(m2_bid),
        .m2_bresp(m2_bresp),
        .m2_bvalid(m2_bvalid),
        .m2_bready(m2_bready),
        .m2_arid(m2_arid),
        .m2_araddr(m2_araddr),
        .m2_arlen(m2_arlen),
        .m2_arsize(m2_arsize),
        .m2_arburst(m2_arburst),
        .m2_arlock(m2_arlock),
        .m2_arcache(m2_arcache),
        .m2_arprot(m2_arprot),
        .m2_arqos(m2_arqos),
        .m2_arvalid(m2_arvalid),
        .m2_arready(m2_arready),
        .m2_rid(m2_rid),
        .m2_rdata(m2_rdata),
        .m2_rresp(m2_rresp),
        .m2_rlast(m2_rlast),
        .m2_rvalid(m2_rvalid),
        .m2_rready(m2_rready),
        // Master 3 connections
        .m3_awid(m3_awid),
        .m3_awaddr(m3_awaddr),
        .m3_awlen(m3_awlen),
        .m3_awsize(m3_awsize),
        .m3_awburst(m3_awburst),
        .m3_awlock(m3_awlock),
        .m3_awcache(m3_awcache),
        .m3_awprot(m3_awprot),
        .m3_awqos(m3_awqos),
        .m3_awvalid(m3_awvalid),
        .m3_awready(m3_awready),
        .m3_wdata(m3_wdata),
        .m3_wstrb(m3_wstrb),
        .m3_wlast(m3_wlast),
        .m3_wvalid(m3_wvalid),
        .m3_wready(m3_wready),
        .m3_bid(m3_bid),
        .m3_bresp(m3_bresp),
        .m3_bvalid(m3_bvalid),
        .m3_bready(m3_bready),
        .m3_arid(m3_arid),
        .m3_araddr(m3_araddr),
        .m3_arlen(m3_arlen),
        .m3_arsize(m3_arsize),
        .m3_arburst(m3_arburst),
        .m3_arlock(m3_arlock),
        .m3_arcache(m3_arcache),
        .m3_arprot(m3_arprot),
        .m3_arqos(m3_arqos),
        .m3_arvalid(m3_arvalid),
        .m3_arready(m3_arready),
        .m3_rid(m3_rid),
        .m3_rdata(m3_rdata),
        .m3_rresp(m3_rresp),
        .m3_rlast(m3_rlast),
        .m3_rvalid(m3_rvalid),
        .m3_rready(m3_rready),
        // Master 4 connections
        .m4_awid(m4_awid),
        .m4_awaddr(m4_awaddr),
        .m4_awlen(m4_awlen),
        .m4_awsize(m4_awsize),
        .m4_awburst(m4_awburst),
        .m4_awlock(m4_awlock),
        .m4_awcache(m4_awcache),
        .m4_awprot(m4_awprot),
        .m4_awqos(m4_awqos),
        .m4_awvalid(m4_awvalid),
        .m4_awready(m4_awready),
        .m4_wdata(m4_wdata),
        .m4_wstrb(m4_wstrb),
        .m4_wlast(m4_wlast),
        .m4_wvalid(m4_wvalid),
        .m4_wready(m4_wready),
        .m4_bid(m4_bid),
        .m4_bresp(m4_bresp),
        .m4_bvalid(m4_bvalid),
        .m4_bready(m4_bready),
        .m4_arid(m4_arid),
        .m4_araddr(m4_araddr),
        .m4_arlen(m4_arlen),
        .m4_arsize(m4_arsize),
        .m4_arburst(m4_arburst),
        .m4_arlock(m4_arlock),
        .m4_arcache(m4_arcache),
        .m4_arprot(m4_arprot),
        .m4_arqos(m4_arqos),
        .m4_arvalid(m4_arvalid),
        .m4_arready(m4_arready),
        .m4_rid(m4_rid),
        .m4_rdata(m4_rdata),
        .m4_rresp(m4_rresp),
        .m4_rlast(m4_rlast),
        .m4_rvalid(m4_rvalid),
        .m4_rready(m4_rready),
        // Master 5 connections
        .m5_awid(m5_awid),
        .m5_awaddr(m5_awaddr),
        .m5_awlen(m5_awlen),
        .m5_awsize(m5_awsize),
        .m5_awburst(m5_awburst),
        .m5_awlock(m5_awlock),
        .m5_awcache(m5_awcache),
        .m5_awprot(m5_awprot),
        .m5_awqos(m5_awqos),
        .m5_awvalid(m5_awvalid),
        .m5_awready(m5_awready),
        .m5_wdata(m5_wdata),
        .m5_wstrb(m5_wstrb),
        .m5_wlast(m5_wlast),
        .m5_wvalid(m5_wvalid),
        .m5_wready(m5_wready),
        .m5_bid(m5_bid),
        .m5_bresp(m5_bresp),
        .m5_bvalid(m5_bvalid),
        .m5_bready(m5_bready),
        .m5_arid(m5_arid),
        .m5_araddr(m5_araddr),
        .m5_arlen(m5_arlen),
        .m5_arsize(m5_arsize),
        .m5_arburst(m5_arburst),
        .m5_arlock(m5_arlock),
        .m5_arcache(m5_arcache),
        .m5_arprot(m5_arprot),
        .m5_arqos(m5_arqos),
        .m5_arvalid(m5_arvalid),
        .m5_arready(m5_arready),
        .m5_rid(m5_rid),
        .m5_rdata(m5_rdata),
        .m5_rresp(m5_rresp),
        .m5_rlast(m5_rlast),
        .m5_rvalid(m5_rvalid),
        .m5_rready(m5_rready),
        // Master 6 connections
        .m6_awid(m6_awid),
        .m6_awaddr(m6_awaddr),
        .m6_awlen(m6_awlen),
        .m6_awsize(m6_awsize),
        .m6_awburst(m6_awburst),
        .m6_awlock(m6_awlock),
        .m6_awcache(m6_awcache),
        .m6_awprot(m6_awprot),
        .m6_awqos(m6_awqos),
        .m6_awvalid(m6_awvalid),
        .m6_awready(m6_awready),
        .m6_wdata(m6_wdata),
        .m6_wstrb(m6_wstrb),
        .m6_wlast(m6_wlast),
        .m6_wvalid(m6_wvalid),
        .m6_wready(m6_wready),
        .m6_bid(m6_bid),
        .m6_bresp(m6_bresp),
        .m6_bvalid(m6_bvalid),
        .m6_bready(m6_bready),
        .m6_arid(m6_arid),
        .m6_araddr(m6_araddr),
        .m6_arlen(m6_arlen),
        .m6_arsize(m6_arsize),
        .m6_arburst(m6_arburst),
        .m6_arlock(m6_arlock),
        .m6_arcache(m6_arcache),
        .m6_arprot(m6_arprot),
        .m6_arqos(m6_arqos),
        .m6_arvalid(m6_arvalid),
        .m6_arready(m6_arready),
        .m6_rid(m6_rid),
        .m6_rdata(m6_rdata),
        .m6_rresp(m6_rresp),
        .m6_rlast(m6_rlast),
        .m6_rvalid(m6_rvalid),
        .m6_rready(m6_rready),
        // Master 7 connections
        .m7_awid(m7_awid),
        .m7_awaddr(m7_awaddr),
        .m7_awlen(m7_awlen),
        .m7_awsize(m7_awsize),
        .m7_awburst(m7_awburst),
        .m7_awlock(m7_awlock),
        .m7_awcache(m7_awcache),
        .m7_awprot(m7_awprot),
        .m7_awqos(m7_awqos),
        .m7_awvalid(m7_awvalid),
        .m7_awready(m7_awready),
        .m7_wdata(m7_wdata),
        .m7_wstrb(m7_wstrb),
        .m7_wlast(m7_wlast),
        .m7_wvalid(m7_wvalid),
        .m7_wready(m7_wready),
        .m7_bid(m7_bid),
        .m7_bresp(m7_bresp),
        .m7_bvalid(m7_bvalid),
        .m7_bready(m7_bready),
        .m7_arid(m7_arid),
        .m7_araddr(m7_araddr),
        .m7_arlen(m7_arlen),
        .m7_arsize(m7_arsize),
        .m7_arburst(m7_arburst),
        .m7_arlock(m7_arlock),
        .m7_arcache(m7_arcache),
        .m7_arprot(m7_arprot),
        .m7_arqos(m7_arqos),
        .m7_arvalid(m7_arvalid),
        .m7_arready(m7_arready),
        .m7_rid(m7_rid),
        .m7_rdata(m7_rdata),
        .m7_rresp(m7_rresp),
        .m7_rlast(m7_rlast),
        .m7_rvalid(m7_rvalid),
        .m7_rready(m7_rready),
        // Master 8 connections
        .m8_awid(m8_awid),
        .m8_awaddr(m8_awaddr),
        .m8_awlen(m8_awlen),
        .m8_awsize(m8_awsize),
        .m8_awburst(m8_awburst),
        .m8_awlock(m8_awlock),
        .m8_awcache(m8_awcache),
        .m8_awprot(m8_awprot),
        .m8_awqos(m8_awqos),
        .m8_awvalid(m8_awvalid),
        .m8_awready(m8_awready),
        .m8_wdata(m8_wdata),
        .m8_wstrb(m8_wstrb),
        .m8_wlast(m8_wlast),
        .m8_wvalid(m8_wvalid),
        .m8_wready(m8_wready),
        .m8_bid(m8_bid),
        .m8_bresp(m8_bresp),
        .m8_bvalid(m8_bvalid),
        .m8_bready(m8_bready),
        .m8_arid(m8_arid),
        .m8_araddr(m8_araddr),
        .m8_arlen(m8_arlen),
        .m8_arsize(m8_arsize),
        .m8_arburst(m8_arburst),
        .m8_arlock(m8_arlock),
        .m8_arcache(m8_arcache),
        .m8_arprot(m8_arprot),
        .m8_arqos(m8_arqos),
        .m8_arvalid(m8_arvalid),
        .m8_arready(m8_arready),
        .m8_rid(m8_rid),
        .m8_rdata(m8_rdata),
        .m8_rresp(m8_rresp),
        .m8_rlast(m8_rlast),
        .m8_rvalid(m8_rvalid),
        .m8_rready(m8_rready),
        // Master 9 connections
        .m9_awid(m9_awid),
        .m9_awaddr(m9_awaddr),
        .m9_awlen(m9_awlen),
        .m9_awsize(m9_awsize),
        .m9_awburst(m9_awburst),
        .m9_awlock(m9_awlock),
        .m9_awcache(m9_awcache),
        .m9_awprot(m9_awprot),
        .m9_awqos(m9_awqos),
        .m9_awvalid(m9_awvalid),
        .m9_awready(m9_awready),
        .m9_wdata(m9_wdata),
        .m9_wstrb(m9_wstrb),
        .m9_wlast(m9_wlast),
        .m9_wvalid(m9_wvalid),
        .m9_wready(m9_wready),
        .m9_bid(m9_bid),
        .m9_bresp(m9_bresp),
        .m9_bvalid(m9_bvalid),
        .m9_bready(m9_bready),
        .m9_arid(m9_arid),
        .m9_araddr(m9_araddr),
        .m9_arlen(m9_arlen),
        .m9_arsize(m9_arsize),
        .m9_arburst(m9_arburst),
        .m9_arlock(m9_arlock),
        .m9_arcache(m9_arcache),
        .m9_arprot(m9_arprot),
        .m9_arqos(m9_arqos),
        .m9_arvalid(m9_arvalid),
        .m9_arready(m9_arready),
        .m9_rid(m9_rid),
        .m9_rdata(m9_rdata),
        .m9_rresp(m9_rresp),
        .m9_rlast(m9_rlast),
        .m9_rvalid(m9_rvalid),
        .m9_rready(m9_rready),
        // Master 10 connections
        .m10_awid(m10_awid),
        .m10_awaddr(m10_awaddr),
        .m10_awlen(m10_awlen),
        .m10_awsize(m10_awsize),
        .m10_awburst(m10_awburst),
        .m10_awlock(m10_awlock),
        .m10_awcache(m10_awcache),
        .m10_awprot(m10_awprot),
        .m10_awqos(m10_awqos),
        .m10_awvalid(m10_awvalid),
        .m10_awready(m10_awready),
        .m10_wdata(m10_wdata),
        .m10_wstrb(m10_wstrb),
        .m10_wlast(m10_wlast),
        .m10_wvalid(m10_wvalid),
        .m10_wready(m10_wready),
        .m10_bid(m10_bid),
        .m10_bresp(m10_bresp),
        .m10_bvalid(m10_bvalid),
        .m10_bready(m10_bready),
        .m10_arid(m10_arid),
        .m10_araddr(m10_araddr),
        .m10_arlen(m10_arlen),
        .m10_arsize(m10_arsize),
        .m10_arburst(m10_arburst),
        .m10_arlock(m10_arlock),
        .m10_arcache(m10_arcache),
        .m10_arprot(m10_arprot),
        .m10_arqos(m10_arqos),
        .m10_arvalid(m10_arvalid),
        .m10_arready(m10_arready),
        .m10_rid(m10_rid),
        .m10_rdata(m10_rdata),
        .m10_rresp(m10_rresp),
        .m10_rlast(m10_rlast),
        .m10_rvalid(m10_rvalid),
        .m10_rready(m10_rready),
        // Master 11 connections
        .m11_awid(m11_awid),
        .m11_awaddr(m11_awaddr),
        .m11_awlen(m11_awlen),
        .m11_awsize(m11_awsize),
        .m11_awburst(m11_awburst),
        .m11_awlock(m11_awlock),
        .m11_awcache(m11_awcache),
        .m11_awprot(m11_awprot),
        .m11_awqos(m11_awqos),
        .m11_awvalid(m11_awvalid),
        .m11_awready(m11_awready),
        .m11_wdata(m11_wdata),
        .m11_wstrb(m11_wstrb),
        .m11_wlast(m11_wlast),
        .m11_wvalid(m11_wvalid),
        .m11_wready(m11_wready),
        .m11_bid(m11_bid),
        .m11_bresp(m11_bresp),
        .m11_bvalid(m11_bvalid),
        .m11_bready(m11_bready),
        .m11_arid(m11_arid),
        .m11_araddr(m11_araddr),
        .m11_arlen(m11_arlen),
        .m11_arsize(m11_arsize),
        .m11_arburst(m11_arburst),
        .m11_arlock(m11_arlock),
        .m11_arcache(m11_arcache),
        .m11_arprot(m11_arprot),
        .m11_arqos(m11_arqos),
        .m11_arvalid(m11_arvalid),
        .m11_arready(m11_arready),
        .m11_rid(m11_rid),
        .m11_rdata(m11_rdata),
        .m11_rresp(m11_rresp),
        .m11_rlast(m11_rlast),
        .m11_rvalid(m11_rvalid),
        .m11_rready(m11_rready),
        // Master 12 connections
        .m12_awid(m12_awid),
        .m12_awaddr(m12_awaddr),
        .m12_awlen(m12_awlen),
        .m12_awsize(m12_awsize),
        .m12_awburst(m12_awburst),
        .m12_awlock(m12_awlock),
        .m12_awcache(m12_awcache),
        .m12_awprot(m12_awprot),
        .m12_awqos(m12_awqos),
        .m12_awvalid(m12_awvalid),
        .m12_awready(m12_awready),
        .m12_wdata(m12_wdata),
        .m12_wstrb(m12_wstrb),
        .m12_wlast(m12_wlast),
        .m12_wvalid(m12_wvalid),
        .m12_wready(m12_wready),
        .m12_bid(m12_bid),
        .m12_bresp(m12_bresp),
        .m12_bvalid(m12_bvalid),
        .m12_bready(m12_bready),
        .m12_arid(m12_arid),
        .m12_araddr(m12_araddr),
        .m12_arlen(m12_arlen),
        .m12_arsize(m12_arsize),
        .m12_arburst(m12_arburst),
        .m12_arlock(m12_arlock),
        .m12_arcache(m12_arcache),
        .m12_arprot(m12_arprot),
        .m12_arqos(m12_arqos),
        .m12_arvalid(m12_arvalid),
        .m12_arready(m12_arready),
        .m12_rid(m12_rid),
        .m12_rdata(m12_rdata),
        .m12_rresp(m12_rresp),
        .m12_rlast(m12_rlast),
        .m12_rvalid(m12_rvalid),
        .m12_rready(m12_rready),
        // Master 13 connections
        .m13_awid(m13_awid),
        .m13_awaddr(m13_awaddr),
        .m13_awlen(m13_awlen),
        .m13_awsize(m13_awsize),
        .m13_awburst(m13_awburst),
        .m13_awlock(m13_awlock),
        .m13_awcache(m13_awcache),
        .m13_awprot(m13_awprot),
        .m13_awqos(m13_awqos),
        .m13_awvalid(m13_awvalid),
        .m13_awready(m13_awready),
        .m13_wdata(m13_wdata),
        .m13_wstrb(m13_wstrb),
        .m13_wlast(m13_wlast),
        .m13_wvalid(m13_wvalid),
        .m13_wready(m13_wready),
        .m13_bid(m13_bid),
        .m13_bresp(m13_bresp),
        .m13_bvalid(m13_bvalid),
        .m13_bready(m13_bready),
        .m13_arid(m13_arid),
        .m13_araddr(m13_araddr),
        .m13_arlen(m13_arlen),
        .m13_arsize(m13_arsize),
        .m13_arburst(m13_arburst),
        .m13_arlock(m13_arlock),
        .m13_arcache(m13_arcache),
        .m13_arprot(m13_arprot),
        .m13_arqos(m13_arqos),
        .m13_arvalid(m13_arvalid),
        .m13_arready(m13_arready),
        .m13_rid(m13_rid),
        .m13_rdata(m13_rdata),
        .m13_rresp(m13_rresp),
        .m13_rlast(m13_rlast),
        .m13_rvalid(m13_rvalid),
        .m13_rready(m13_rready),
        // Master 14 connections
        .m14_awid(m14_awid),
        .m14_awaddr(m14_awaddr),
        .m14_awlen(m14_awlen),
        .m14_awsize(m14_awsize),
        .m14_awburst(m14_awburst),
        .m14_awlock(m14_awlock),
        .m14_awcache(m14_awcache),
        .m14_awprot(m14_awprot),
        .m14_awqos(m14_awqos),
        .m14_awvalid(m14_awvalid),
        .m14_awready(m14_awready),
        .m14_wdata(m14_wdata),
        .m14_wstrb(m14_wstrb),
        .m14_wlast(m14_wlast),
        .m14_wvalid(m14_wvalid),
        .m14_wready(m14_wready),
        .m14_bid(m14_bid),
        .m14_bresp(m14_bresp),
        .m14_bvalid(m14_bvalid),
        .m14_bready(m14_bready),
        .m14_arid(m14_arid),
        .m14_araddr(m14_araddr),
        .m14_arlen(m14_arlen),
        .m14_arsize(m14_arsize),
        .m14_arburst(m14_arburst),
        .m14_arlock(m14_arlock),
        .m14_arcache(m14_arcache),
        .m14_arprot(m14_arprot),
        .m14_arqos(m14_arqos),
        .m14_arvalid(m14_arvalid),
        .m14_arready(m14_arready),
        .m14_rid(m14_rid),
        .m14_rdata(m14_rdata),
        .m14_rresp(m14_rresp),
        .m14_rlast(m14_rlast),
        .m14_rvalid(m14_rvalid),
        .m14_rready(m14_rready),
        // Slave 0 connections
        .s0_awid(s0_awid),
        .s0_awaddr(s0_awaddr),
        .s0_awlen(s0_awlen),
        .s0_awsize(s0_awsize),
        .s0_awburst(s0_awburst),
        .s0_awlock(s0_awlock),
        .s0_awcache(s0_awcache),
        .s0_awprot(s0_awprot),
        .s0_awqos(s0_awqos),
        .s0_awvalid(s0_awvalid),
        .s0_awready(s0_awready),
        .s0_wdata(s0_wdata),
        .s0_wstrb(s0_wstrb),
        .s0_wlast(s0_wlast),
        .s0_wvalid(s0_wvalid),
        .s0_wready(s0_wready),
        .s0_bid(s0_bid),
        .s0_bresp(s0_bresp),
        .s0_bvalid(s0_bvalid),
        .s0_bready(s0_bready),
        .s0_arid(s0_arid),
        .s0_araddr(s0_araddr),
        .s0_arlen(s0_arlen),
        .s0_arsize(s0_arsize),
        .s0_arburst(s0_arburst),
        .s0_arlock(s0_arlock),
        .s0_arcache(s0_arcache),
        .s0_arprot(s0_arprot),
        .s0_arqos(s0_arqos),
        .s0_arvalid(s0_arvalid),
        .s0_arready(s0_arready),
        .s0_rid(s0_rid),
        .s0_rdata(s0_rdata),
        .s0_rresp(s0_rresp),
        .s0_rlast(s0_rlast),
        .s0_rvalid(s0_rvalid),
        .s0_rready(s0_rready),
        // Slave 1 connections
        .s1_awid(s1_awid),
        .s1_awaddr(s1_awaddr),
        .s1_awlen(s1_awlen),
        .s1_awsize(s1_awsize),
        .s1_awburst(s1_awburst),
        .s1_awlock(s1_awlock),
        .s1_awcache(s1_awcache),
        .s1_awprot(s1_awprot),
        .s1_awqos(s1_awqos),
        .s1_awvalid(s1_awvalid),
        .s1_awready(s1_awready),
        .s1_wdata(s1_wdata),
        .s1_wstrb(s1_wstrb),
        .s1_wlast(s1_wlast),
        .s1_wvalid(s1_wvalid),
        .s1_wready(s1_wready),
        .s1_bid(s1_bid),
        .s1_bresp(s1_bresp),
        .s1_bvalid(s1_bvalid),
        .s1_bready(s1_bready),
        .s1_arid(s1_arid),
        .s1_araddr(s1_araddr),
        .s1_arlen(s1_arlen),
        .s1_arsize(s1_arsize),
        .s1_arburst(s1_arburst),
        .s1_arlock(s1_arlock),
        .s1_arcache(s1_arcache),
        .s1_arprot(s1_arprot),
        .s1_arqos(s1_arqos),
        .s1_arvalid(s1_arvalid),
        .s1_arready(s1_arready),
        .s1_rid(s1_rid),
        .s1_rdata(s1_rdata),
        .s1_rresp(s1_rresp),
        .s1_rlast(s1_rlast),
        .s1_rvalid(s1_rvalid),
        .s1_rready(s1_rready),
        // Slave 2 connections
        .s2_awid(s2_awid),
        .s2_awaddr(s2_awaddr),
        .s2_awlen(s2_awlen),
        .s2_awsize(s2_awsize),
        .s2_awburst(s2_awburst),
        .s2_awlock(s2_awlock),
        .s2_awcache(s2_awcache),
        .s2_awprot(s2_awprot),
        .s2_awqos(s2_awqos),
        .s2_awvalid(s2_awvalid),
        .s2_awready(s2_awready),
        .s2_wdata(s2_wdata),
        .s2_wstrb(s2_wstrb),
        .s2_wlast(s2_wlast),
        .s2_wvalid(s2_wvalid),
        .s2_wready(s2_wready),
        .s2_bid(s2_bid),
        .s2_bresp(s2_bresp),
        .s2_bvalid(s2_bvalid),
        .s2_bready(s2_bready),
        .s2_arid(s2_arid),
        .s2_araddr(s2_araddr),
        .s2_arlen(s2_arlen),
        .s2_arsize(s2_arsize),
        .s2_arburst(s2_arburst),
        .s2_arlock(s2_arlock),
        .s2_arcache(s2_arcache),
        .s2_arprot(s2_arprot),
        .s2_arqos(s2_arqos),
        .s2_arvalid(s2_arvalid),
        .s2_arready(s2_arready),
        .s2_rid(s2_rid),
        .s2_rdata(s2_rdata),
        .s2_rresp(s2_rresp),
        .s2_rlast(s2_rlast),
        .s2_rvalid(s2_rvalid),
        .s2_rready(s2_rready),
        // Slave 3 connections
        .s3_awid(s3_awid),
        .s3_awaddr(s3_awaddr),
        .s3_awlen(s3_awlen),
        .s3_awsize(s3_awsize),
        .s3_awburst(s3_awburst),
        .s3_awlock(s3_awlock),
        .s3_awcache(s3_awcache),
        .s3_awprot(s3_awprot),
        .s3_awqos(s3_awqos),
        .s3_awvalid(s3_awvalid),
        .s3_awready(s3_awready),
        .s3_wdata(s3_wdata),
        .s3_wstrb(s3_wstrb),
        .s3_wlast(s3_wlast),
        .s3_wvalid(s3_wvalid),
        .s3_wready(s3_wready),
        .s3_bid(s3_bid),
        .s3_bresp(s3_bresp),
        .s3_bvalid(s3_bvalid),
        .s3_bready(s3_bready),
        .s3_arid(s3_arid),
        .s3_araddr(s3_araddr),
        .s3_arlen(s3_arlen),
        .s3_arsize(s3_arsize),
        .s3_arburst(s3_arburst),
        .s3_arlock(s3_arlock),
        .s3_arcache(s3_arcache),
        .s3_arprot(s3_arprot),
        .s3_arqos(s3_arqos),
        .s3_arvalid(s3_arvalid),
        .s3_arready(s3_arready),
        .s3_rid(s3_rid),
        .s3_rdata(s3_rdata),
        .s3_rresp(s3_rresp),
        .s3_rlast(s3_rlast),
        .s3_rvalid(s3_rvalid),
        .s3_rready(s3_rready),
        // Slave 4 connections
        .s4_awid(s4_awid),
        .s4_awaddr(s4_awaddr),
        .s4_awlen(s4_awlen),
        .s4_awsize(s4_awsize),
        .s4_awburst(s4_awburst),
        .s4_awlock(s4_awlock),
        .s4_awcache(s4_awcache),
        .s4_awprot(s4_awprot),
        .s4_awqos(s4_awqos),
        .s4_awvalid(s4_awvalid),
        .s4_awready(s4_awready),
        .s4_wdata(s4_wdata),
        .s4_wstrb(s4_wstrb),
        .s4_wlast(s4_wlast),
        .s4_wvalid(s4_wvalid),
        .s4_wready(s4_wready),
        .s4_bid(s4_bid),
        .s4_bresp(s4_bresp),
        .s4_bvalid(s4_bvalid),
        .s4_bready(s4_bready),
        .s4_arid(s4_arid),
        .s4_araddr(s4_araddr),
        .s4_arlen(s4_arlen),
        .s4_arsize(s4_arsize),
        .s4_arburst(s4_arburst),
        .s4_arlock(s4_arlock),
        .s4_arcache(s4_arcache),
        .s4_arprot(s4_arprot),
        .s4_arqos(s4_arqos),
        .s4_arvalid(s4_arvalid),
        .s4_arready(s4_arready),
        .s4_rid(s4_rid),
        .s4_rdata(s4_rdata),
        .s4_rresp(s4_rresp),
        .s4_rlast(s4_rlast),
        .s4_rvalid(s4_rvalid),
        .s4_rready(s4_rready),
        // Slave 5 connections
        .s5_awid(s5_awid),
        .s5_awaddr(s5_awaddr),
        .s5_awlen(s5_awlen),
        .s5_awsize(s5_awsize),
        .s5_awburst(s5_awburst),
        .s5_awlock(s5_awlock),
        .s5_awcache(s5_awcache),
        .s5_awprot(s5_awprot),
        .s5_awqos(s5_awqos),
        .s5_awvalid(s5_awvalid),
        .s5_awready(s5_awready),
        .s5_wdata(s5_wdata),
        .s5_wstrb(s5_wstrb),
        .s5_wlast(s5_wlast),
        .s5_wvalid(s5_wvalid),
        .s5_wready(s5_wready),
        .s5_bid(s5_bid),
        .s5_bresp(s5_bresp),
        .s5_bvalid(s5_bvalid),
        .s5_bready(s5_bready),
        .s5_arid(s5_arid),
        .s5_araddr(s5_araddr),
        .s5_arlen(s5_arlen),
        .s5_arsize(s5_arsize),
        .s5_arburst(s5_arburst),
        .s5_arlock(s5_arlock),
        .s5_arcache(s5_arcache),
        .s5_arprot(s5_arprot),
        .s5_arqos(s5_arqos),
        .s5_arvalid(s5_arvalid),
        .s5_arready(s5_arready),
        .s5_rid(s5_rid),
        .s5_rdata(s5_rdata),
        .s5_rresp(s5_rresp),
        .s5_rlast(s5_rlast),
        .s5_rvalid(s5_rvalid),
        .s5_rready(s5_rready),
        // Slave 6 connections
        .s6_awid(s6_awid),
        .s6_awaddr(s6_awaddr),
        .s6_awlen(s6_awlen),
        .s6_awsize(s6_awsize),
        .s6_awburst(s6_awburst),
        .s6_awlock(s6_awlock),
        .s6_awcache(s6_awcache),
        .s6_awprot(s6_awprot),
        .s6_awqos(s6_awqos),
        .s6_awvalid(s6_awvalid),
        .s6_awready(s6_awready),
        .s6_wdata(s6_wdata),
        .s6_wstrb(s6_wstrb),
        .s6_wlast(s6_wlast),
        .s6_wvalid(s6_wvalid),
        .s6_wready(s6_wready),
        .s6_bid(s6_bid),
        .s6_bresp(s6_bresp),
        .s6_bvalid(s6_bvalid),
        .s6_bready(s6_bready),
        .s6_arid(s6_arid),
        .s6_araddr(s6_araddr),
        .s6_arlen(s6_arlen),
        .s6_arsize(s6_arsize),
        .s6_arburst(s6_arburst),
        .s6_arlock(s6_arlock),
        .s6_arcache(s6_arcache),
        .s6_arprot(s6_arprot),
        .s6_arqos(s6_arqos),
        .s6_arvalid(s6_arvalid),
        .s6_arready(s6_arready),
        .s6_rid(s6_rid),
        .s6_rdata(s6_rdata),
        .s6_rresp(s6_rresp),
        .s6_rlast(s6_rlast),
        .s6_rvalid(s6_rvalid),
        .s6_rready(s6_rready),
        // Slave 7 connections
        .s7_awid(s7_awid),
        .s7_awaddr(s7_awaddr),
        .s7_awlen(s7_awlen),
        .s7_awsize(s7_awsize),
        .s7_awburst(s7_awburst),
        .s7_awlock(s7_awlock),
        .s7_awcache(s7_awcache),
        .s7_awprot(s7_awprot),
        .s7_awqos(s7_awqos),
        .s7_awvalid(s7_awvalid),
        .s7_awready(s7_awready),
        .s7_wdata(s7_wdata),
        .s7_wstrb(s7_wstrb),
        .s7_wlast(s7_wlast),
        .s7_wvalid(s7_wvalid),
        .s7_wready(s7_wready),
        .s7_bid(s7_bid),
        .s7_bresp(s7_bresp),
        .s7_bvalid(s7_bvalid),
        .s7_bready(s7_bready),
        .s7_arid(s7_arid),
        .s7_araddr(s7_araddr),
        .s7_arlen(s7_arlen),
        .s7_arsize(s7_arsize),
        .s7_arburst(s7_arburst),
        .s7_arlock(s7_arlock),
        .s7_arcache(s7_arcache),
        .s7_arprot(s7_arprot),
        .s7_arqos(s7_arqos),
        .s7_arvalid(s7_arvalid),
        .s7_arready(s7_arready),
        .s7_rid(s7_rid),
        .s7_rdata(s7_rdata),
        .s7_rresp(s7_rresp),
        .s7_rlast(s7_rlast),
        .s7_rvalid(s7_rvalid),
        .s7_rready(s7_rready),
        // Slave 8 connections
        .s8_awid(s8_awid),
        .s8_awaddr(s8_awaddr),
        .s8_awlen(s8_awlen),
        .s8_awsize(s8_awsize),
        .s8_awburst(s8_awburst),
        .s8_awlock(s8_awlock),
        .s8_awcache(s8_awcache),
        .s8_awprot(s8_awprot),
        .s8_awqos(s8_awqos),
        .s8_awvalid(s8_awvalid),
        .s8_awready(s8_awready),
        .s8_wdata(s8_wdata),
        .s8_wstrb(s8_wstrb),
        .s8_wlast(s8_wlast),
        .s8_wvalid(s8_wvalid),
        .s8_wready(s8_wready),
        .s8_bid(s8_bid),
        .s8_bresp(s8_bresp),
        .s8_bvalid(s8_bvalid),
        .s8_bready(s8_bready),
        .s8_arid(s8_arid),
        .s8_araddr(s8_araddr),
        .s8_arlen(s8_arlen),
        .s8_arsize(s8_arsize),
        .s8_arburst(s8_arburst),
        .s8_arlock(s8_arlock),
        .s8_arcache(s8_arcache),
        .s8_arprot(s8_arprot),
        .s8_arqos(s8_arqos),
        .s8_arvalid(s8_arvalid),
        .s8_arready(s8_arready),
        .s8_rid(s8_rid),
        .s8_rdata(s8_rdata),
        .s8_rresp(s8_rresp),
        .s8_rlast(s8_rlast),
        .s8_rvalid(s8_rvalid),
        .s8_rready(s8_rready),
        // Slave 9 connections
        .s9_awid(s9_awid),
        .s9_awaddr(s9_awaddr),
        .s9_awlen(s9_awlen),
        .s9_awsize(s9_awsize),
        .s9_awburst(s9_awburst),
        .s9_awlock(s9_awlock),
        .s9_awcache(s9_awcache),
        .s9_awprot(s9_awprot),
        .s9_awqos(s9_awqos),
        .s9_awvalid(s9_awvalid),
        .s9_awready(s9_awready),
        .s9_wdata(s9_wdata),
        .s9_wstrb(s9_wstrb),
        .s9_wlast(s9_wlast),
        .s9_wvalid(s9_wvalid),
        .s9_wready(s9_wready),
        .s9_bid(s9_bid),
        .s9_bresp(s9_bresp),
        .s9_bvalid(s9_bvalid),
        .s9_bready(s9_bready),
        .s9_arid(s9_arid),
        .s9_araddr(s9_araddr),
        .s9_arlen(s9_arlen),
        .s9_arsize(s9_arsize),
        .s9_arburst(s9_arburst),
        .s9_arlock(s9_arlock),
        .s9_arcache(s9_arcache),
        .s9_arprot(s9_arprot),
        .s9_arqos(s9_arqos),
        .s9_arvalid(s9_arvalid),
        .s9_arready(s9_arready),
        .s9_rid(s9_rid),
        .s9_rdata(s9_rdata),
        .s9_rresp(s9_rresp),
        .s9_rlast(s9_rlast),
        .s9_rvalid(s9_rvalid),
        .s9_rready(s9_rready),
        // Slave 10 connections
        .s10_awid(s10_awid),
        .s10_awaddr(s10_awaddr),
        .s10_awlen(s10_awlen),
        .s10_awsize(s10_awsize),
        .s10_awburst(s10_awburst),
        .s10_awlock(s10_awlock),
        .s10_awcache(s10_awcache),
        .s10_awprot(s10_awprot),
        .s10_awqos(s10_awqos),
        .s10_awvalid(s10_awvalid),
        .s10_awready(s10_awready),
        .s10_wdata(s10_wdata),
        .s10_wstrb(s10_wstrb),
        .s10_wlast(s10_wlast),
        .s10_wvalid(s10_wvalid),
        .s10_wready(s10_wready),
        .s10_bid(s10_bid),
        .s10_bresp(s10_bresp),
        .s10_bvalid(s10_bvalid),
        .s10_bready(s10_bready),
        .s10_arid(s10_arid),
        .s10_araddr(s10_araddr),
        .s10_arlen(s10_arlen),
        .s10_arsize(s10_arsize),
        .s10_arburst(s10_arburst),
        .s10_arlock(s10_arlock),
        .s10_arcache(s10_arcache),
        .s10_arprot(s10_arprot),
        .s10_arqos(s10_arqos),
        .s10_arvalid(s10_arvalid),
        .s10_arready(s10_arready),
        .s10_rid(s10_rid),
        .s10_rdata(s10_rdata),
        .s10_rresp(s10_rresp),
        .s10_rlast(s10_rlast),
        .s10_rvalid(s10_rvalid),
        .s10_rready(s10_rready),
        // Slave 11 connections
        .s11_awid(s11_awid),
        .s11_awaddr(s11_awaddr),
        .s11_awlen(s11_awlen),
        .s11_awsize(s11_awsize),
        .s11_awburst(s11_awburst),
        .s11_awlock(s11_awlock),
        .s11_awcache(s11_awcache),
        .s11_awprot(s11_awprot),
        .s11_awqos(s11_awqos),
        .s11_awvalid(s11_awvalid),
        .s11_awready(s11_awready),
        .s11_wdata(s11_wdata),
        .s11_wstrb(s11_wstrb),
        .s11_wlast(s11_wlast),
        .s11_wvalid(s11_wvalid),
        .s11_wready(s11_wready),
        .s11_bid(s11_bid),
        .s11_bresp(s11_bresp),
        .s11_bvalid(s11_bvalid),
        .s11_bready(s11_bready),
        .s11_arid(s11_arid),
        .s11_araddr(s11_araddr),
        .s11_arlen(s11_arlen),
        .s11_arsize(s11_arsize),
        .s11_arburst(s11_arburst),
        .s11_arlock(s11_arlock),
        .s11_arcache(s11_arcache),
        .s11_arprot(s11_arprot),
        .s11_arqos(s11_arqos),
        .s11_arvalid(s11_arvalid),
        .s11_arready(s11_arready),
        .s11_rid(s11_rid),
        .s11_rdata(s11_rdata),
        .s11_rresp(s11_rresp),
        .s11_rlast(s11_rlast),
        .s11_rvalid(s11_rvalid),
        .s11_rready(s11_rready),
        // Slave 12 connections
        .s12_awid(s12_awid),
        .s12_awaddr(s12_awaddr),
        .s12_awlen(s12_awlen),
        .s12_awsize(s12_awsize),
        .s12_awburst(s12_awburst),
        .s12_awlock(s12_awlock),
        .s12_awcache(s12_awcache),
        .s12_awprot(s12_awprot),
        .s12_awqos(s12_awqos),
        .s12_awvalid(s12_awvalid),
        .s12_awready(s12_awready),
        .s12_wdata(s12_wdata),
        .s12_wstrb(s12_wstrb),
        .s12_wlast(s12_wlast),
        .s12_wvalid(s12_wvalid),
        .s12_wready(s12_wready),
        .s12_bid(s12_bid),
        .s12_bresp(s12_bresp),
        .s12_bvalid(s12_bvalid),
        .s12_bready(s12_bready),
        .s12_arid(s12_arid),
        .s12_araddr(s12_araddr),
        .s12_arlen(s12_arlen),
        .s12_arsize(s12_arsize),
        .s12_arburst(s12_arburst),
        .s12_arlock(s12_arlock),
        .s12_arcache(s12_arcache),
        .s12_arprot(s12_arprot),
        .s12_arqos(s12_arqos),
        .s12_arvalid(s12_arvalid),
        .s12_arready(s12_arready),
        .s12_rid(s12_rid),
        .s12_rdata(s12_rdata),
        .s12_rresp(s12_rresp),
        .s12_rlast(s12_rlast),
        .s12_rvalid(s12_rvalid),
        .s12_rready(s12_rready),
        // Slave 13 connections
        .s13_awid(s13_awid),
        .s13_awaddr(s13_awaddr),
        .s13_awlen(s13_awlen),
        .s13_awsize(s13_awsize),
        .s13_awburst(s13_awburst),
        .s13_awlock(s13_awlock),
        .s13_awcache(s13_awcache),
        .s13_awprot(s13_awprot),
        .s13_awqos(s13_awqos),
        .s13_awvalid(s13_awvalid),
        .s13_awready(s13_awready),
        .s13_wdata(s13_wdata),
        .s13_wstrb(s13_wstrb),
        .s13_wlast(s13_wlast),
        .s13_wvalid(s13_wvalid),
        .s13_wready(s13_wready),
        .s13_bid(s13_bid),
        .s13_bresp(s13_bresp),
        .s13_bvalid(s13_bvalid),
        .s13_bready(s13_bready),
        .s13_arid(s13_arid),
        .s13_araddr(s13_araddr),
        .s13_arlen(s13_arlen),
        .s13_arsize(s13_arsize),
        .s13_arburst(s13_arburst),
        .s13_arlock(s13_arlock),
        .s13_arcache(s13_arcache),
        .s13_arprot(s13_arprot),
        .s13_arqos(s13_arqos),
        .s13_arvalid(s13_arvalid),
        .s13_arready(s13_arready),
        .s13_rid(s13_rid),
        .s13_rdata(s13_rdata),
        .s13_rresp(s13_rresp),
        .s13_rlast(s13_rlast),
        .s13_rvalid(s13_rvalid),
        .s13_rready(s13_rready),
        // Slave 14 connections
        .s14_awid(s14_awid),
        .s14_awaddr(s14_awaddr),
        .s14_awlen(s14_awlen),
        .s14_awsize(s14_awsize),
        .s14_awburst(s14_awburst),
        .s14_awlock(s14_awlock),
        .s14_awcache(s14_awcache),
        .s14_awprot(s14_awprot),
        .s14_awqos(s14_awqos),
        .s14_awvalid(s14_awvalid),
        .s14_awready(s14_awready),
        .s14_wdata(s14_wdata),
        .s14_wstrb(s14_wstrb),
        .s14_wlast(s14_wlast),
        .s14_wvalid(s14_wvalid),
        .s14_wready(s14_wready),
        .s14_bid(s14_bid),
        .s14_bresp(s14_bresp),
        .s14_bvalid(s14_bvalid),
        .s14_bready(s14_bready),
        .s14_arid(s14_arid),
        .s14_araddr(s14_araddr),
        .s14_arlen(s14_arlen),
        .s14_arsize(s14_arsize),
        .s14_arburst(s14_arburst),
        .s14_arlock(s14_arlock),
        .s14_arcache(s14_arcache),
        .s14_arprot(s14_arprot),
        .s14_arqos(s14_arqos),
        .s14_arvalid(s14_arvalid),
        .s14_arready(s14_arready),
        .s14_rid(s14_rid),
        .s14_rdata(s14_rdata),
        .s14_rresp(s14_rresp),
        .s14_rlast(s14_rlast),
        .s14_rvalid(s14_rvalid),
        .s14_rready(s14_rready)
