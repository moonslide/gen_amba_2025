// Wrapper module to adapt between VIP and gen_amba_axi naming conventions
// This wrapper translates signal names from the VIP testbench format
// to the format expected by the generated RTL

module axi4_interconnect_m9s9 #(
    parameter DATA_WIDTH = 64,
    parameter ADDR_WIDTH = 32,
    parameter ID_WIDTH = 4
)(
    // Clock and reset - VIP format
    input  logic                      aclk,
    input  logic                      aresetn,
    
    // Master 0 AXI interface - VIP format
    input  logic [ID_WIDTH-1:0]       m0_awid,
    input  logic [ADDR_WIDTH-1:0]     m0_awaddr,
    input  logic [7:0]                m0_awlen,
    input  logic [2:0]                m0_awsize,
    input  logic [1:0]                m0_awburst,
    input  logic                      m0_awlock,
    input  logic [3:0]                m0_awcache,
    input  logic [2:0]                m0_awprot,
    input  logic [3:0]                m0_awqos,
    input  logic                      m0_awvalid,
    output logic                      m0_awready,
    
    input  logic [DATA_WIDTH-1:0]     m0_wdata,
    input  logic [DATA_WIDTH/8-1:0]   m0_wstrb,
    input  logic                      m0_wlast,
    input  logic                      m0_wvalid,
    output logic                      m0_wready,
    
    output logic [ID_WIDTH-1:0]       m0_bid,
    output logic [1:0]                m0_bresp,
    output logic                      m0_bvalid,
    input  logic                      m0_bready,
    
    input  logic [ID_WIDTH-1:0]       m0_arid,
    input  logic [ADDR_WIDTH-1:0]     m0_araddr,
    input  logic [7:0]                m0_arlen,
    input  logic [2:0]                m0_arsize,
    input  logic [1:0]                m0_arburst,
    input  logic                      m0_arlock,
    input  logic [3:0]                m0_arcache,
    input  logic [2:0]                m0_arprot,
    input  logic [3:0]                m0_arqos,
    input  logic                      m0_arvalid,
    output logic                      m0_arready,
    
    output logic [ID_WIDTH-1:0]       m0_rid,
    output logic [DATA_WIDTH-1:0]     m0_rdata,
    output logic [1:0]                m0_rresp,
    output logic                      m0_rlast,
    output logic                      m0_rvalid,
    input  logic                      m0_rready,
    
    // Master 1 interface
    input  logic [ID_WIDTH-1:0]       m1_awid,
    input  logic [ADDR_WIDTH-1:0]     m1_awaddr,
    input  logic [7:0]                m1_awlen,
    input  logic [2:0]                m1_awsize,
    input  logic [1:0]                m1_awburst,
    input  logic                      m1_awlock,
    input  logic [3:0]                m1_awcache,
    input  logic [2:0]                m1_awprot,
    input  logic [3:0]                m1_awqos,
    input  logic                      m1_awvalid,
    output logic                      m1_awready,
    input  logic [DATA_WIDTH-1:0]     m1_wdata,
    input  logic [DATA_WIDTH/8-1:0]   m1_wstrb,
    input  logic                      m1_wlast,
    input  logic                      m1_wvalid,
    output logic                      m1_wready,
    output logic [ID_WIDTH-1:0]       m1_bid,
    output logic [1:0]                m1_bresp,
    output logic                      m1_bvalid,
    input  logic                      m1_bready,
    input  logic [ID_WIDTH-1:0]       m1_arid,
    input  logic [ADDR_WIDTH-1:0]     m1_araddr,
    input  logic [7:0]                m1_arlen,
    input  logic [2:0]                m1_arsize,
    input  logic [1:0]                m1_arburst,
    input  logic                      m1_arlock,
    input  logic [3:0]                m1_arcache,
    input  logic [2:0]                m1_arprot,
    input  logic [3:0]                m1_arqos,
    input  logic                      m1_arvalid,
    output logic                      m1_arready,
    output logic [ID_WIDTH-1:0]       m1_rid,
    output logic [DATA_WIDTH-1:0]     m1_rdata,
    output logic [1:0]                m1_rresp,
    output logic                      m1_rlast,
    output logic                      m1_rvalid,
    input  logic                      m1_rready,
    
    // Master 2-8 interfaces (abbreviated for space - same pattern)
    // M2
    input  logic [ID_WIDTH-1:0]       m2_awid,
    input  logic [ADDR_WIDTH-1:0]     m2_awaddr,
    input  logic [7:0]                m2_awlen,
    input  logic [2:0]                m2_awsize,
    input  logic [1:0]                m2_awburst,
    input  logic                      m2_awlock,
    input  logic [3:0]                m2_awcache,
    input  logic [2:0]                m2_awprot,
    input  logic [3:0]                m2_awqos,
    input  logic                      m2_awvalid,
    output logic                      m2_awready,
    input  logic [DATA_WIDTH-1:0]     m2_wdata,
    input  logic [DATA_WIDTH/8-1:0]   m2_wstrb,
    input  logic                      m2_wlast,
    input  logic                      m2_wvalid,
    output logic                      m2_wready,
    output logic [ID_WIDTH-1:0]       m2_bid,
    output logic [1:0]                m2_bresp,
    output logic                      m2_bvalid,
    input  logic                      m2_bready,
    input  logic [ID_WIDTH-1:0]       m2_arid,
    input  logic [ADDR_WIDTH-1:0]     m2_araddr,
    input  logic [7:0]                m2_arlen,
    input  logic [2:0]                m2_arsize,
    input  logic [1:0]                m2_arburst,
    input  logic                      m2_arlock,
    input  logic [3:0]                m2_arcache,
    input  logic [2:0]                m2_arprot,
    input  logic [3:0]                m2_arqos,
    input  logic                      m2_arvalid,
    output logic                      m2_arready,
    output logic [ID_WIDTH-1:0]       m2_rid,
    output logic [DATA_WIDTH-1:0]     m2_rdata,
    output logic [1:0]                m2_rresp,
    output logic                      m2_rlast,
    output logic                      m2_rvalid,
    input  logic                      m2_rready,
    
    // M3
    input  logic [ID_WIDTH-1:0]       m3_awid,
    input  logic [ADDR_WIDTH-1:0]     m3_awaddr,
    input  logic [7:0]                m3_awlen,
    input  logic [2:0]                m3_awsize,
    input  logic [1:0]                m3_awburst,
    input  logic                      m3_awlock,
    input  logic [3:0]                m3_awcache,
    input  logic [2:0]                m3_awprot,
    input  logic [3:0]                m3_awqos,
    input  logic                      m3_awvalid,
    output logic                      m3_awready,
    input  logic [DATA_WIDTH-1:0]     m3_wdata,
    input  logic [DATA_WIDTH/8-1:0]   m3_wstrb,
    input  logic                      m3_wlast,
    input  logic                      m3_wvalid,
    output logic                      m3_wready,
    output logic [ID_WIDTH-1:0]       m3_bid,
    output logic [1:0]                m3_bresp,
    output logic                      m3_bvalid,
    input  logic                      m3_bready,
    input  logic [ID_WIDTH-1:0]       m3_arid,
    input  logic [ADDR_WIDTH-1:0]     m3_araddr,
    input  logic [7:0]                m3_arlen,
    input  logic [2:0]                m3_arsize,
    input  logic [1:0]                m3_arburst,
    input  logic                      m3_arlock,
    input  logic [3:0]                m3_arcache,
    input  logic [2:0]                m3_arprot,
    input  logic [3:0]                m3_arqos,
    input  logic                      m3_arvalid,
    output logic                      m3_arready,
    output logic [ID_WIDTH-1:0]       m3_rid,
    output logic [DATA_WIDTH-1:0]     m3_rdata,
    output logic [1:0]                m3_rresp,
    output logic                      m3_rlast,
    output logic                      m3_rvalid,
    input  logic                      m3_rready,
    
    // M4
    input  logic [ID_WIDTH-1:0]       m4_awid,
    input  logic [ADDR_WIDTH-1:0]     m4_awaddr,
    input  logic [7:0]                m4_awlen,
    input  logic [2:0]                m4_awsize,
    input  logic [1:0]                m4_awburst,
    input  logic                      m4_awlock,
    input  logic [3:0]                m4_awcache,
    input  logic [2:0]                m4_awprot,
    input  logic [3:0]                m4_awqos,
    input  logic                      m4_awvalid,
    output logic                      m4_awready,
    input  logic [DATA_WIDTH-1:0]     m4_wdata,
    input  logic [DATA_WIDTH/8-1:0]   m4_wstrb,
    input  logic                      m4_wlast,
    input  logic                      m4_wvalid,
    output logic                      m4_wready,
    output logic [ID_WIDTH-1:0]       m4_bid,
    output logic [1:0]                m4_bresp,
    output logic                      m4_bvalid,
    input  logic                      m4_bready,
    input  logic [ID_WIDTH-1:0]       m4_arid,
    input  logic [ADDR_WIDTH-1:0]     m4_araddr,
    input  logic [7:0]                m4_arlen,
    input  logic [2:0]                m4_arsize,
    input  logic [1:0]                m4_arburst,
    input  logic                      m4_arlock,
    input  logic [3:0]                m4_arcache,
    input  logic [2:0]                m4_arprot,
    input  logic [3:0]                m4_arqos,
    input  logic                      m4_arvalid,
    output logic                      m4_arready,
    output logic [ID_WIDTH-1:0]       m4_rid,
    output logic [DATA_WIDTH-1:0]     m4_rdata,
    output logic [1:0]                m4_rresp,
    output logic                      m4_rlast,
    output logic                      m4_rvalid,
    input  logic                      m4_rready,
    
    // M5
    input  logic [ID_WIDTH-1:0]       m5_awid,
    input  logic [ADDR_WIDTH-1:0]     m5_awaddr,
    input  logic [7:0]                m5_awlen,
    input  logic [2:0]                m5_awsize,
    input  logic [1:0]                m5_awburst,
    input  logic                      m5_awlock,
    input  logic [3:0]                m5_awcache,
    input  logic [2:0]                m5_awprot,
    input  logic [3:0]                m5_awqos,
    input  logic                      m5_awvalid,
    output logic                      m5_awready,
    input  logic [DATA_WIDTH-1:0]     m5_wdata,
    input  logic [DATA_WIDTH/8-1:0]   m5_wstrb,
    input  logic                      m5_wlast,
    input  logic                      m5_wvalid,
    output logic                      m5_wready,
    output logic [ID_WIDTH-1:0]       m5_bid,
    output logic [1:0]                m5_bresp,
    output logic                      m5_bvalid,
    input  logic                      m5_bready,
    input  logic [ID_WIDTH-1:0]       m5_arid,
    input  logic [ADDR_WIDTH-1:0]     m5_araddr,
    input  logic [7:0]                m5_arlen,
    input  logic [2:0]                m5_arsize,
    input  logic [1:0]                m5_arburst,
    input  logic                      m5_arlock,
    input  logic [3:0]                m5_arcache,
    input  logic [2:0]                m5_arprot,
    input  logic [3:0]                m5_arqos,
    input  logic                      m5_arvalid,
    output logic                      m5_arready,
    output logic [ID_WIDTH-1:0]       m5_rid,
    output logic [DATA_WIDTH-1:0]     m5_rdata,
    output logic [1:0]                m5_rresp,
    output logic                      m5_rlast,
    output logic                      m5_rvalid,
    input  logic                      m5_rready,
    
    // M6
    input  logic [ID_WIDTH-1:0]       m6_awid,
    input  logic [ADDR_WIDTH-1:0]     m6_awaddr,
    input  logic [7:0]                m6_awlen,
    input  logic [2:0]                m6_awsize,
    input  logic [1:0]                m6_awburst,
    input  logic                      m6_awlock,
    input  logic [3:0]                m6_awcache,
    input  logic [2:0]                m6_awprot,
    input  logic [3:0]                m6_awqos,
    input  logic                      m6_awvalid,
    output logic                      m6_awready,
    input  logic [DATA_WIDTH-1:0]     m6_wdata,
    input  logic [DATA_WIDTH/8-1:0]   m6_wstrb,
    input  logic                      m6_wlast,
    input  logic                      m6_wvalid,
    output logic                      m6_wready,
    output logic [ID_WIDTH-1:0]       m6_bid,
    output logic [1:0]                m6_bresp,
    output logic                      m6_bvalid,
    input  logic                      m6_bready,
    input  logic [ID_WIDTH-1:0]       m6_arid,
    input  logic [ADDR_WIDTH-1:0]     m6_araddr,
    input  logic [7:0]                m6_arlen,
    input  logic [2:0]                m6_arsize,
    input  logic [1:0]                m6_arburst,
    input  logic                      m6_arlock,
    input  logic [3:0]                m6_arcache,
    input  logic [2:0]                m6_arprot,
    input  logic [3:0]                m6_arqos,
    input  logic                      m6_arvalid,
    output logic                      m6_arready,
    output logic [ID_WIDTH-1:0]       m6_rid,
    output logic [DATA_WIDTH-1:0]     m6_rdata,
    output logic [1:0]                m6_rresp,
    output logic                      m6_rlast,
    output logic                      m6_rvalid,
    input  logic                      m6_rready,
    
    // M7
    input  logic [ID_WIDTH-1:0]       m7_awid,
    input  logic [ADDR_WIDTH-1:0]     m7_awaddr,
    input  logic [7:0]                m7_awlen,
    input  logic [2:0]                m7_awsize,
    input  logic [1:0]                m7_awburst,
    input  logic                      m7_awlock,
    input  logic [3:0]                m7_awcache,
    input  logic [2:0]                m7_awprot,
    input  logic [3:0]                m7_awqos,
    input  logic                      m7_awvalid,
    output logic                      m7_awready,
    input  logic [DATA_WIDTH-1:0]     m7_wdata,
    input  logic [DATA_WIDTH/8-1:0]   m7_wstrb,
    input  logic                      m7_wlast,
    input  logic                      m7_wvalid,
    output logic                      m7_wready,
    output logic [ID_WIDTH-1:0]       m7_bid,
    output logic [1:0]                m7_bresp,
    output logic                      m7_bvalid,
    input  logic                      m7_bready,
    input  logic [ID_WIDTH-1:0]       m7_arid,
    input  logic [ADDR_WIDTH-1:0]     m7_araddr,
    input  logic [7:0]                m7_arlen,
    input  logic [2:0]                m7_arsize,
    input  logic [1:0]                m7_arburst,
    input  logic                      m7_arlock,
    input  logic [3:0]                m7_arcache,
    input  logic [2:0]                m7_arprot,
    input  logic [3:0]                m7_arqos,
    input  logic                      m7_arvalid,
    output logic                      m7_arready,
    output logic [ID_WIDTH-1:0]       m7_rid,
    output logic [DATA_WIDTH-1:0]     m7_rdata,
    output logic [1:0]                m7_rresp,
    output logic                      m7_rlast,
    output logic                      m7_rvalid,
    input  logic                      m7_rready,
    
    // M8
    input  logic [ID_WIDTH-1:0]       m8_awid,
    input  logic [ADDR_WIDTH-1:0]     m8_awaddr,
    input  logic [7:0]                m8_awlen,
    input  logic [2:0]                m8_awsize,
    input  logic [1:0]                m8_awburst,
    input  logic                      m8_awlock,
    input  logic [3:0]                m8_awcache,
    input  logic [2:0]                m8_awprot,
    input  logic [3:0]                m8_awqos,
    input  logic                      m8_awvalid,
    output logic                      m8_awready,
    input  logic [DATA_WIDTH-1:0]     m8_wdata,
    input  logic [DATA_WIDTH/8-1:0]   m8_wstrb,
    input  logic                      m8_wlast,
    input  logic                      m8_wvalid,
    output logic                      m8_wready,
    output logic [ID_WIDTH-1:0]       m8_bid,
    output logic [1:0]                m8_bresp,
    output logic                      m8_bvalid,
    input  logic                      m8_bready,
    input  logic [ID_WIDTH-1:0]       m8_arid,
    input  logic [ADDR_WIDTH-1:0]     m8_araddr,
    input  logic [7:0]                m8_arlen,
    input  logic [2:0]                m8_arsize,
    input  logic [1:0]                m8_arburst,
    input  logic                      m8_arlock,
    input  logic [3:0]                m8_arcache,
    input  logic [2:0]                m8_arprot,
    input  logic [3:0]                m8_arqos,
    input  logic                      m8_arvalid,
    output logic                      m8_arready,
    output logic [ID_WIDTH-1:0]       m8_rid,
    output logic [DATA_WIDTH-1:0]     m8_rdata,
    output logic [1:0]                m8_rresp,
    output logic                      m8_rlast,
    output logic                      m8_rvalid,
    input  logic                      m8_rready,
    
    // Slave 0 AXI interface - VIP format
    output logic [ID_WIDTH+$clog2(9)-1:0] s0_awid,
    output logic [ADDR_WIDTH-1:0]     s0_awaddr,
    output logic [7:0]                s0_awlen,
    output logic [2:0]                s0_awsize,
    output logic [1:0]                s0_awburst,
    output logic                      s0_awlock,
    output logic [3:0]                s0_awcache,
    output logic [2:0]                s0_awprot,
    output logic [3:0]                s0_awqos,
    output logic                      s0_awvalid,
    input  logic                      s0_awready,
    
    output logic [DATA_WIDTH-1:0]     s0_wdata,
    output logic [DATA_WIDTH/8-1:0]   s0_wstrb,
    output logic                      s0_wlast,
    output logic                      s0_wvalid,
    input  logic                      s0_wready,
    
    input  logic [ID_WIDTH+$clog2(9)-1:0] s0_bid,
    input  logic [1:0]                s0_bresp,
    input  logic                      s0_bvalid,
    output logic                      s0_bready,
    
    output logic [ID_WIDTH+$clog2(9)-1:0] s0_arid,
    output logic [ADDR_WIDTH-1:0]     s0_araddr,
    output logic [7:0]                s0_arlen,
    output logic [2:0]                s0_arsize,
    output logic [1:0]                s0_arburst,
    output logic                      s0_arlock,
    output logic [3:0]                s0_arcache,
    output logic [2:0]                s0_arprot,
    output logic [3:0]                s0_arqos,
    output logic                      s0_arvalid,
    input  logic                      s0_arready,
    
    input  logic [ID_WIDTH+$clog2(9)-1:0] s0_rid,
    input  logic [DATA_WIDTH-1:0]     s0_rdata,
    input  logic [1:0]                s0_rresp,
    input  logic                      s0_rlast,
    input  logic                      s0_rvalid,
    output logic                      s0_rready,
    
    // Slave 1-8 (same pattern)
    // S1
    output logic [ID_WIDTH+$clog2(9)-1:0] s1_awid,
    output logic [ADDR_WIDTH-1:0]     s1_awaddr,
    output logic [7:0]                s1_awlen,
    output logic [2:0]                s1_awsize,
    output logic [1:0]                s1_awburst,
    output logic                      s1_awlock,
    output logic [3:0]                s1_awcache,
    output logic [2:0]                s1_awprot,
    output logic [3:0]                s1_awqos,
    output logic                      s1_awvalid,
    input  logic                      s1_awready,
    output logic [DATA_WIDTH-1:0]     s1_wdata,
    output logic [DATA_WIDTH/8-1:0]   s1_wstrb,
    output logic                      s1_wlast,
    output logic                      s1_wvalid,
    input  logic                      s1_wready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s1_bid,
    input  logic [1:0]                s1_bresp,
    input  logic                      s1_bvalid,
    output logic                      s1_bready,
    output logic [ID_WIDTH+$clog2(9)-1:0] s1_arid,
    output logic [ADDR_WIDTH-1:0]     s1_araddr,
    output logic [7:0]                s1_arlen,
    output logic [2:0]                s1_arsize,
    output logic [1:0]                s1_arburst,
    output logic                      s1_arlock,
    output logic [3:0]                s1_arcache,
    output logic [2:0]                s1_arprot,
    output logic [3:0]                s1_arqos,
    output logic                      s1_arvalid,
    input  logic                      s1_arready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s1_rid,
    input  logic [DATA_WIDTH-1:0]     s1_rdata,
    input  logic [1:0]                s1_rresp,
    input  logic                      s1_rlast,
    input  logic                      s1_rvalid,
    output logic                      s1_rready,
    
    // S2
    output logic [ID_WIDTH+$clog2(9)-1:0] s2_awid,
    output logic [ADDR_WIDTH-1:0]     s2_awaddr,
    output logic [7:0]                s2_awlen,
    output logic [2:0]                s2_awsize,
    output logic [1:0]                s2_awburst,
    output logic                      s2_awlock,
    output logic [3:0]                s2_awcache,
    output logic [2:0]                s2_awprot,
    output logic [3:0]                s2_awqos,
    output logic                      s2_awvalid,
    input  logic                      s2_awready,
    output logic [DATA_WIDTH-1:0]     s2_wdata,
    output logic [DATA_WIDTH/8-1:0]   s2_wstrb,
    output logic                      s2_wlast,
    output logic                      s2_wvalid,
    input  logic                      s2_wready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s2_bid,
    input  logic [1:0]                s2_bresp,
    input  logic                      s2_bvalid,
    output logic                      s2_bready,
    output logic [ID_WIDTH+$clog2(9)-1:0] s2_arid,
    output logic [ADDR_WIDTH-1:0]     s2_araddr,
    output logic [7:0]                s2_arlen,
    output logic [2:0]                s2_arsize,
    output logic [1:0]                s2_arburst,
    output logic                      s2_arlock,
    output logic [3:0]                s2_arcache,
    output logic [2:0]                s2_arprot,
    output logic [3:0]                s2_arqos,
    output logic                      s2_arvalid,
    input  logic                      s2_arready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s2_rid,
    input  logic [DATA_WIDTH-1:0]     s2_rdata,
    input  logic [1:0]                s2_rresp,
    input  logic                      s2_rlast,
    input  logic                      s2_rvalid,
    output logic                      s2_rready,
    
    // S3
    output logic [ID_WIDTH+$clog2(9)-1:0] s3_awid,
    output logic [ADDR_WIDTH-1:0]     s3_awaddr,
    output logic [7:0]                s3_awlen,
    output logic [2:0]                s3_awsize,
    output logic [1:0]                s3_awburst,
    output logic                      s3_awlock,
    output logic [3:0]                s3_awcache,
    output logic [2:0]                s3_awprot,
    output logic [3:0]                s3_awqos,
    output logic                      s3_awvalid,
    input  logic                      s3_awready,
    output logic [DATA_WIDTH-1:0]     s3_wdata,
    output logic [DATA_WIDTH/8-1:0]   s3_wstrb,
    output logic                      s3_wlast,
    output logic                      s3_wvalid,
    input  logic                      s3_wready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s3_bid,
    input  logic [1:0]                s3_bresp,
    input  logic                      s3_bvalid,
    output logic                      s3_bready,
    output logic [ID_WIDTH+$clog2(9)-1:0] s3_arid,
    output logic [ADDR_WIDTH-1:0]     s3_araddr,
    output logic [7:0]                s3_arlen,
    output logic [2:0]                s3_arsize,
    output logic [1:0]                s3_arburst,
    output logic                      s3_arlock,
    output logic [3:0]                s3_arcache,
    output logic [2:0]                s3_arprot,
    output logic [3:0]                s3_arqos,
    output logic                      s3_arvalid,
    input  logic                      s3_arready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s3_rid,
    input  logic [DATA_WIDTH-1:0]     s3_rdata,
    input  logic [1:0]                s3_rresp,
    input  logic                      s3_rlast,
    input  logic                      s3_rvalid,
    output logic                      s3_rready,
    
    // S4
    output logic [ID_WIDTH+$clog2(9)-1:0] s4_awid,
    output logic [ADDR_WIDTH-1:0]     s4_awaddr,
    output logic [7:0]                s4_awlen,
    output logic [2:0]                s4_awsize,
    output logic [1:0]                s4_awburst,
    output logic                      s4_awlock,
    output logic [3:0]                s4_awcache,
    output logic [2:0]                s4_awprot,
    output logic [3:0]                s4_awqos,
    output logic                      s4_awvalid,
    input  logic                      s4_awready,
    output logic [DATA_WIDTH-1:0]     s4_wdata,
    output logic [DATA_WIDTH/8-1:0]   s4_wstrb,
    output logic                      s4_wlast,
    output logic                      s4_wvalid,
    input  logic                      s4_wready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s4_bid,
    input  logic [1:0]                s4_bresp,
    input  logic                      s4_bvalid,
    output logic                      s4_bready,
    output logic [ID_WIDTH+$clog2(9)-1:0] s4_arid,
    output logic [ADDR_WIDTH-1:0]     s4_araddr,
    output logic [7:0]                s4_arlen,
    output logic [2:0]                s4_arsize,
    output logic [1:0]                s4_arburst,
    output logic                      s4_arlock,
    output logic [3:0]                s4_arcache,
    output logic [2:0]                s4_arprot,
    output logic [3:0]                s4_arqos,
    output logic                      s4_arvalid,
    input  logic                      s4_arready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s4_rid,
    input  logic [DATA_WIDTH-1:0]     s4_rdata,
    input  logic [1:0]                s4_rresp,
    input  logic                      s4_rlast,
    input  logic                      s4_rvalid,
    output logic                      s4_rready,
    
    // S5
    output logic [ID_WIDTH+$clog2(9)-1:0] s5_awid,
    output logic [ADDR_WIDTH-1:0]     s5_awaddr,
    output logic [7:0]                s5_awlen,
    output logic [2:0]                s5_awsize,
    output logic [1:0]                s5_awburst,
    output logic                      s5_awlock,
    output logic [3:0]                s5_awcache,
    output logic [2:0]                s5_awprot,
    output logic [3:0]                s5_awqos,
    output logic                      s5_awvalid,
    input  logic                      s5_awready,
    output logic [DATA_WIDTH-1:0]     s5_wdata,
    output logic [DATA_WIDTH/8-1:0]   s5_wstrb,
    output logic                      s5_wlast,
    output logic                      s5_wvalid,
    input  logic                      s5_wready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s5_bid,
    input  logic [1:0]                s5_bresp,
    input  logic                      s5_bvalid,
    output logic                      s5_bready,
    output logic [ID_WIDTH+$clog2(9)-1:0] s5_arid,
    output logic [ADDR_WIDTH-1:0]     s5_araddr,
    output logic [7:0]                s5_arlen,
    output logic [2:0]                s5_arsize,
    output logic [1:0]                s5_arburst,
    output logic                      s5_arlock,
    output logic [3:0]                s5_arcache,
    output logic [2:0]                s5_arprot,
    output logic [3:0]                s5_arqos,
    output logic                      s5_arvalid,
    input  logic                      s5_arready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s5_rid,
    input  logic [DATA_WIDTH-1:0]     s5_rdata,
    input  logic [1:0]                s5_rresp,
    input  logic                      s5_rlast,
    input  logic                      s5_rvalid,
    output logic                      s5_rready,
    
    // S6
    output logic [ID_WIDTH+$clog2(9)-1:0] s6_awid,
    output logic [ADDR_WIDTH-1:0]     s6_awaddr,
    output logic [7:0]                s6_awlen,
    output logic [2:0]                s6_awsize,
    output logic [1:0]                s6_awburst,
    output logic                      s6_awlock,
    output logic [3:0]                s6_awcache,
    output logic [2:0]                s6_awprot,
    output logic [3:0]                s6_awqos,
    output logic                      s6_awvalid,
    input  logic                      s6_awready,
    output logic [DATA_WIDTH-1:0]     s6_wdata,
    output logic [DATA_WIDTH/8-1:0]   s6_wstrb,
    output logic                      s6_wlast,
    output logic                      s6_wvalid,
    input  logic                      s6_wready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s6_bid,
    input  logic [1:0]                s6_bresp,
    input  logic                      s6_bvalid,
    output logic                      s6_bready,
    output logic [ID_WIDTH+$clog2(9)-1:0] s6_arid,
    output logic [ADDR_WIDTH-1:0]     s6_araddr,
    output logic [7:0]                s6_arlen,
    output logic [2:0]                s6_arsize,
    output logic [1:0]                s6_arburst,
    output logic                      s6_arlock,
    output logic [3:0]                s6_arcache,
    output logic [2:0]                s6_arprot,
    output logic [3:0]                s6_arqos,
    output logic                      s6_arvalid,
    input  logic                      s6_arready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s6_rid,
    input  logic [DATA_WIDTH-1:0]     s6_rdata,
    input  logic [1:0]                s6_rresp,
    input  logic                      s6_rlast,
    input  logic                      s6_rvalid,
    output logic                      s6_rready,
    
    // S7
    output logic [ID_WIDTH+$clog2(9)-1:0] s7_awid,
    output logic [ADDR_WIDTH-1:0]     s7_awaddr,
    output logic [7:0]                s7_awlen,
    output logic [2:0]                s7_awsize,
    output logic [1:0]                s7_awburst,
    output logic                      s7_awlock,
    output logic [3:0]                s7_awcache,
    output logic [2:0]                s7_awprot,
    output logic [3:0]                s7_awqos,
    output logic                      s7_awvalid,
    input  logic                      s7_awready,
    output logic [DATA_WIDTH-1:0]     s7_wdata,
    output logic [DATA_WIDTH/8-1:0]   s7_wstrb,
    output logic                      s7_wlast,
    output logic                      s7_wvalid,
    input  logic                      s7_wready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s7_bid,
    input  logic [1:0]                s7_bresp,
    input  logic                      s7_bvalid,
    output logic                      s7_bready,
    output logic [ID_WIDTH+$clog2(9)-1:0] s7_arid,
    output logic [ADDR_WIDTH-1:0]     s7_araddr,
    output logic [7:0]                s7_arlen,
    output logic [2:0]                s7_arsize,
    output logic [1:0]                s7_arburst,
    output logic                      s7_arlock,
    output logic [3:0]                s7_arcache,
    output logic [2:0]                s7_arprot,
    output logic [3:0]                s7_arqos,
    output logic                      s7_arvalid,
    input  logic                      s7_arready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s7_rid,
    input  logic [DATA_WIDTH-1:0]     s7_rdata,
    input  logic [1:0]                s7_rresp,
    input  logic                      s7_rlast,
    input  logic                      s7_rvalid,
    output logic                      s7_rready,
    
    // S8
    output logic [ID_WIDTH+$clog2(9)-1:0] s8_awid,
    output logic [ADDR_WIDTH-1:0]     s8_awaddr,
    output logic [7:0]                s8_awlen,
    output logic [2:0]                s8_awsize,
    output logic [1:0]                s8_awburst,
    output logic                      s8_awlock,
    output logic [3:0]                s8_awcache,
    output logic [2:0]                s8_awprot,
    output logic [3:0]                s8_awqos,
    output logic                      s8_awvalid,
    input  logic                      s8_awready,
    output logic [DATA_WIDTH-1:0]     s8_wdata,
    output logic [DATA_WIDTH/8-1:0]   s8_wstrb,
    output logic                      s8_wlast,
    output logic                      s8_wvalid,
    input  logic                      s8_wready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s8_bid,
    input  logic [1:0]                s8_bresp,
    input  logic                      s8_bvalid,
    output logic                      s8_bready,
    output logic [ID_WIDTH+$clog2(9)-1:0] s8_arid,
    output logic [ADDR_WIDTH-1:0]     s8_araddr,
    output logic [7:0]                s8_arlen,
    output logic [2:0]                s8_arsize,
    output logic [1:0]                s8_arburst,
    output logic                      s8_arlock,
    output logic [3:0]                s8_arcache,
    output logic [2:0]                s8_arprot,
    output logic [3:0]                s8_arqos,
    output logic                      s8_arvalid,
    input  logic                      s8_arready,
    input  logic [ID_WIDTH+$clog2(9)-1:0] s8_rid,
    input  logic [DATA_WIDTH-1:0]     s8_rdata,
    input  logic [1:0]                s8_rresp,
    input  logic                      s8_rlast,
    input  logic                      s8_rvalid,
    output logic                      s8_rready
);

    // Define macros for conditional compilation
    `define AMBA_AXI_CACHE
    `define AMBA_AXI_PROT
    `define AMBA_QOS
    
    // Instantiate the actual gen_amba_axi interconnect
    amba_axi_m9s9 #(
        .NUM_MASTER  (9),
        .NUM_SLAVE   (9),
        .WIDTH_CID   ($clog2(9)),
        .WIDTH_ID    (ID_WIDTH),
        .WIDTH_AD    (ADDR_WIDTH),
        .WIDTH_DA    (DATA_WIDTH),
        .WIDTH_DS    (DATA_WIDTH/8),
        .WIDTH_SID   ($clog2(9)+ID_WIDTH),
        // Enable all slaves with 4KB address space each
        .SLAVE_EN0(1), .ADDR_LENGTH0(12),
        .SLAVE_EN1(1), .ADDR_LENGTH1(12),
        .SLAVE_EN2(1), .ADDR_LENGTH2(12),
        .SLAVE_EN3(1), .ADDR_LENGTH3(12),
        .SLAVE_EN4(1), .ADDR_LENGTH4(12),
        .SLAVE_EN5(1), .ADDR_LENGTH5(12),
        .SLAVE_EN6(1), .ADDR_LENGTH6(12),
        .SLAVE_EN7(1), .ADDR_LENGTH7(12),
        .SLAVE_EN8(1), .ADDR_LENGTH8(12),
        // Base addresses
        .ADDR_BASE0(32'h00000000),
        .ADDR_BASE1(32'h00001000),
        .ADDR_BASE2(32'h00002000),
        .ADDR_BASE3(32'h00003000),
        .ADDR_BASE4(32'h00004000),
        .ADDR_BASE5(32'h00005000),
        .ADDR_BASE6(32'h00006000),
        .ADDR_BASE7(32'h00007000),
        .ADDR_BASE8(32'h00008000)
    ) u_interconnect (
        // Clock and reset - map naming
        .ARESETn     (aresetn),
        .ACLK        (aclk),
        
        // Master 0 - map all signals
        .M0_AWID     (m0_awid),
        .M0_AWADDR   (m0_awaddr),
        .M0_AWLEN    (m0_awlen),
        .M0_AWSIZE   (m0_awsize),
        .M0_AWBURST  (m0_awburst),
        .M0_AWLOCK   (m0_awlock),
        .M0_AWCACHE  (m0_awcache),
        .M0_AWPROT   (m0_awprot),
        .M0_AWQOS    (m0_awqos),
        .M0_AWREGION (4'b0000),  // Default region
        .M0_AWVALID  (m0_awvalid),
        .M0_AWREADY  (m0_awready),
        .M0_WDATA    (m0_wdata),
        .M0_WSTRB    (m0_wstrb),
        .M0_WLAST    (m0_wlast),
        .M0_WVALID   (m0_wvalid),
        .M0_WREADY   (m0_wready),
        .M0_BID      (m0_bid),
        .M0_BRESP    (m0_bresp),
        .M0_BVALID   (m0_bvalid),
        .M0_BREADY   (m0_bready),
        .M0_ARID     (m0_arid),
        .M0_ARADDR   (m0_araddr),
        .M0_ARLEN    (m0_arlen),
        .M0_ARSIZE   (m0_arsize),
        .M0_ARBURST  (m0_arburst),
        .M0_ARLOCK   (m0_arlock),
        .M0_ARCACHE  (m0_arcache),
        .M0_ARPROT   (m0_arprot),
        .M0_ARQOS    (m0_arqos),
        .M0_ARREGION (4'b0000),
        .M0_ARVALID  (m0_arvalid),
        .M0_ARREADY  (m0_arready),
        .M0_RID      (m0_rid),
        .M0_RDATA    (m0_rdata),
        .M0_RRESP    (m0_rresp),
        .M0_RLAST    (m0_rlast),
        .M0_RVALID   (m0_rvalid),
        .M0_RREADY   (m0_rready),
        
        // Master 1
        .M1_AWID     (m1_awid),
        .M1_AWADDR   (m1_awaddr),
        .M1_AWLEN    (m1_awlen),
        .M1_AWSIZE   (m1_awsize),
        .M1_AWBURST  (m1_awburst),
        .M1_AWLOCK   (m1_awlock),
        .M1_AWCACHE  (m1_awcache),
        .M1_AWPROT   (m1_awprot),
        .M1_AWQOS    (m1_awqos),
        .M1_AWREGION (4'b0000),
        .M1_AWVALID  (m1_awvalid),
        .M1_AWREADY  (m1_awready),
        .M1_WDATA    (m1_wdata),
        .M1_WSTRB    (m1_wstrb),
        .M1_WLAST    (m1_wlast),
        .M1_WVALID   (m1_wvalid),
        .M1_WREADY   (m1_wready),
        .M1_BID      (m1_bid),
        .M1_BRESP    (m1_bresp),
        .M1_BVALID   (m1_bvalid),
        .M1_BREADY   (m1_bready),
        .M1_ARID     (m1_arid),
        .M1_ARADDR   (m1_araddr),
        .M1_ARLEN    (m1_arlen),
        .M1_ARSIZE   (m1_arsize),
        .M1_ARBURST  (m1_arburst),
        .M1_ARLOCK   (m1_arlock),
        .M1_ARCACHE  (m1_arcache),
        .M1_ARPROT   (m1_arprot),
        .M1_ARQOS    (m1_arqos),
        .M1_ARREGION (4'b0000),
        .M1_ARVALID  (m1_arvalid),
        .M1_ARREADY  (m1_arready),
        .M1_RID      (m1_rid),
        .M1_RDATA    (m1_rdata),
        .M1_RRESP    (m1_rresp),
        .M1_RLAST    (m1_rlast),
        .M1_RVALID   (m1_rvalid),
        .M1_RREADY   (m1_rready),
        
        // Master 2
        .M2_AWID     (m2_awid),
        .M2_AWADDR   (m2_awaddr),
        .M2_AWLEN    (m2_awlen),
        .M2_AWSIZE   (m2_awsize),
        .M2_AWBURST  (m2_awburst),
        .M2_AWLOCK   (m2_awlock),
        .M2_AWCACHE  (m2_awcache),
        .M2_AWPROT   (m2_awprot),
        .M2_AWQOS    (m2_awqos),
        .M2_AWREGION (4'b0000),
        .M2_AWVALID  (m2_awvalid),
        .M2_AWREADY  (m2_awready),
        .M2_WDATA    (m2_wdata),
        .M2_WSTRB    (m2_wstrb),
        .M2_WLAST    (m2_wlast),
        .M2_WVALID   (m2_wvalid),
        .M2_WREADY   (m2_wready),
        .M2_BID      (m2_bid),
        .M2_BRESP    (m2_bresp),
        .M2_BVALID   (m2_bvalid),
        .M2_BREADY   (m2_bready),
        .M2_ARID     (m2_arid),
        .M2_ARADDR   (m2_araddr),
        .M2_ARLEN    (m2_arlen),
        .M2_ARSIZE   (m2_arsize),
        .M2_ARBURST  (m2_arburst),
        .M2_ARLOCK   (m2_arlock),
        .M2_ARCACHE  (m2_arcache),
        .M2_ARPROT   (m2_arprot),
        .M2_ARQOS    (m2_arqos),
        .M2_ARREGION (4'b0000),
        .M2_ARVALID  (m2_arvalid),
        .M2_ARREADY  (m2_arready),
        .M2_RID      (m2_rid),
        .M2_RDATA    (m2_rdata),
        .M2_RRESP    (m2_rresp),
        .M2_RLAST    (m2_rlast),
        .M2_RVALID   (m2_rvalid),
        .M2_RREADY   (m2_rready),
        
        // Master 3
        .M3_AWID     (m3_awid),
        .M3_AWADDR   (m3_awaddr),
        .M3_AWLEN    (m3_awlen),
        .M3_AWSIZE   (m3_awsize),
        .M3_AWBURST  (m3_awburst),
        .M3_AWLOCK   (m3_awlock),
        .M3_AWCACHE  (m3_awcache),
        .M3_AWPROT   (m3_awprot),
        .M3_AWQOS    (m3_awqos),
        .M3_AWREGION (4'b0000),
        .M3_AWVALID  (m3_awvalid),
        .M3_AWREADY  (m3_awready),
        .M3_WDATA    (m3_wdata),
        .M3_WSTRB    (m3_wstrb),
        .M3_WLAST    (m3_wlast),
        .M3_WVALID   (m3_wvalid),
        .M3_WREADY   (m3_wready),
        .M3_BID      (m3_bid),
        .M3_BRESP    (m3_bresp),
        .M3_BVALID   (m3_bvalid),
        .M3_BREADY   (m3_bready),
        .M3_ARID     (m3_arid),
        .M3_ARADDR   (m3_araddr),
        .M3_ARLEN    (m3_arlen),
        .M3_ARSIZE   (m3_arsize),
        .M3_ARBURST  (m3_arburst),
        .M3_ARLOCK   (m3_arlock),
        .M3_ARCACHE  (m3_arcache),
        .M3_ARPROT   (m3_arprot),
        .M3_ARQOS    (m3_arqos),
        .M3_ARREGION (4'b0000),
        .M3_ARVALID  (m3_arvalid),
        .M3_ARREADY  (m3_arready),
        .M3_RID      (m3_rid),
        .M3_RDATA    (m3_rdata),
        .M3_RRESP    (m3_rresp),
        .M3_RLAST    (m3_rlast),
        .M3_RVALID   (m3_rvalid),
        .M3_RREADY   (m3_rready),
        
        // Master 4
        .M4_AWID     (m4_awid),
        .M4_AWADDR   (m4_awaddr),
        .M4_AWLEN    (m4_awlen),
        .M4_AWSIZE   (m4_awsize),
        .M4_AWBURST  (m4_awburst),
        .M4_AWLOCK   (m4_awlock),
        .M4_AWCACHE  (m4_awcache),
        .M4_AWPROT   (m4_awprot),
        .M4_AWQOS    (m4_awqos),
        .M4_AWREGION (4'b0000),
        .M4_AWVALID  (m4_awvalid),
        .M4_AWREADY  (m4_awready),
        .M4_WDATA    (m4_wdata),
        .M4_WSTRB    (m4_wstrb),
        .M4_WLAST    (m4_wlast),
        .M4_WVALID   (m4_wvalid),
        .M4_WREADY   (m4_wready),
        .M4_BID      (m4_bid),
        .M4_BRESP    (m4_bresp),
        .M4_BVALID   (m4_bvalid),
        .M4_BREADY   (m4_bready),
        .M4_ARID     (m4_arid),
        .M4_ARADDR   (m4_araddr),
        .M4_ARLEN    (m4_arlen),
        .M4_ARSIZE   (m4_arsize),
        .M4_ARBURST  (m4_arburst),
        .M4_ARLOCK   (m4_arlock),
        .M4_ARCACHE  (m4_arcache),
        .M4_ARPROT   (m4_arprot),
        .M4_ARQOS    (m4_arqos),
        .M4_ARREGION (4'b0000),
        .M4_ARVALID  (m4_arvalid),
        .M4_ARREADY  (m4_arready),
        .M4_RID      (m4_rid),
        .M4_RDATA    (m4_rdata),
        .M4_RRESP    (m4_rresp),
        .M4_RLAST    (m4_rlast),
        .M4_RVALID   (m4_rvalid),
        .M4_RREADY   (m4_rready),
        
        // Master 5
        .M5_AWID     (m5_awid),
        .M5_AWADDR   (m5_awaddr),
        .M5_AWLEN    (m5_awlen),
        .M5_AWSIZE   (m5_awsize),
        .M5_AWBURST  (m5_awburst),
        .M5_AWLOCK   (m5_awlock),
        .M5_AWCACHE  (m5_awcache),
        .M5_AWPROT   (m5_awprot),
        .M5_AWQOS    (m5_awqos),
        .M5_AWREGION (4'b0000),
        .M5_AWVALID  (m5_awvalid),
        .M5_AWREADY  (m5_awready),
        .M5_WDATA    (m5_wdata),
        .M5_WSTRB    (m5_wstrb),
        .M5_WLAST    (m5_wlast),
        .M5_WVALID   (m5_wvalid),
        .M5_WREADY   (m5_wready),
        .M5_BID      (m5_bid),
        .M5_BRESP    (m5_bresp),
        .M5_BVALID   (m5_bvalid),
        .M5_BREADY   (m5_bready),
        .M5_ARID     (m5_arid),
        .M5_ARADDR   (m5_araddr),
        .M5_ARLEN    (m5_arlen),
        .M5_ARSIZE   (m5_arsize),
        .M5_ARBURST  (m5_arburst),
        .M5_ARLOCK   (m5_arlock),
        .M5_ARCACHE  (m5_arcache),
        .M5_ARPROT   (m5_arprot),
        .M5_ARQOS    (m5_arqos),
        .M5_ARREGION (4'b0000),
        .M5_ARVALID  (m5_arvalid),
        .M5_ARREADY  (m5_arready),
        .M5_RID      (m5_rid),
        .M5_RDATA    (m5_rdata),
        .M5_RRESP    (m5_rresp),
        .M5_RLAST    (m5_rlast),
        .M5_RVALID   (m5_rvalid),
        .M5_RREADY   (m5_rready),
        
        // Master 6
        .M6_AWID     (m6_awid),
        .M6_AWADDR   (m6_awaddr),
        .M6_AWLEN    (m6_awlen),
        .M6_AWSIZE   (m6_awsize),
        .M6_AWBURST  (m6_awburst),
        .M6_AWLOCK   (m6_awlock),
        .M6_AWCACHE  (m6_awcache),
        .M6_AWPROT   (m6_awprot),
        .M6_AWQOS    (m6_awqos),
        .M6_AWREGION (4'b0000),
        .M6_AWVALID  (m6_awvalid),
        .M6_AWREADY  (m6_awready),
        .M6_WDATA    (m6_wdata),
        .M6_WSTRB    (m6_wstrb),
        .M6_WLAST    (m6_wlast),
        .M6_WVALID   (m6_wvalid),
        .M6_WREADY   (m6_wready),
        .M6_BID      (m6_bid),
        .M6_BRESP    (m6_bresp),
        .M6_BVALID   (m6_bvalid),
        .M6_BREADY   (m6_bready),
        .M6_ARID     (m6_arid),
        .M6_ARADDR   (m6_araddr),
        .M6_ARLEN    (m6_arlen),
        .M6_ARSIZE   (m6_arsize),
        .M6_ARBURST  (m6_arburst),
        .M6_ARLOCK   (m6_arlock),
        .M6_ARCACHE  (m6_arcache),
        .M6_ARPROT   (m6_arprot),
        .M6_ARQOS    (m6_arqos),
        .M6_ARREGION (4'b0000),
        .M6_ARVALID  (m6_arvalid),
        .M6_ARREADY  (m6_arready),
        .M6_RID      (m6_rid),
        .M6_RDATA    (m6_rdata),
        .M6_RRESP    (m6_rresp),
        .M6_RLAST    (m6_rlast),
        .M6_RVALID   (m6_rvalid),
        .M6_RREADY   (m6_rready),
        
        // Master 7
        .M7_AWID     (m7_awid),
        .M7_AWADDR   (m7_awaddr),
        .M7_AWLEN    (m7_awlen),
        .M7_AWSIZE   (m7_awsize),
        .M7_AWBURST  (m7_awburst),
        .M7_AWLOCK   (m7_awlock),
        .M7_AWCACHE  (m7_awcache),
        .M7_AWPROT   (m7_awprot),
        .M7_AWQOS    (m7_awqos),
        .M7_AWREGION (4'b0000),
        .M7_AWVALID  (m7_awvalid),
        .M7_AWREADY  (m7_awready),
        .M7_WDATA    (m7_wdata),
        .M7_WSTRB    (m7_wstrb),
        .M7_WLAST    (m7_wlast),
        .M7_WVALID   (m7_wvalid),
        .M7_WREADY   (m7_wready),
        .M7_BID      (m7_bid),
        .M7_BRESP    (m7_bresp),
        .M7_BVALID   (m7_bvalid),
        .M7_BREADY   (m7_bready),
        .M7_ARID     (m7_arid),
        .M7_ARADDR   (m7_araddr),
        .M7_ARLEN    (m7_arlen),
        .M7_ARSIZE   (m7_arsize),
        .M7_ARBURST  (m7_arburst),
        .M7_ARLOCK   (m7_arlock),
        .M7_ARCACHE  (m7_arcache),
        .M7_ARPROT   (m7_arprot),
        .M7_ARQOS    (m7_arqos),
        .M7_ARREGION (4'b0000),
        .M7_ARVALID  (m7_arvalid),
        .M7_ARREADY  (m7_arready),
        .M7_RID      (m7_rid),
        .M7_RDATA    (m7_rdata),
        .M7_RRESP    (m7_rresp),
        .M7_RLAST    (m7_rlast),
        .M7_RVALID   (m7_rvalid),
        .M7_RREADY   (m7_rready),
        
        // Master 8
        .M8_AWID     (m8_awid),
        .M8_AWADDR   (m8_awaddr),
        .M8_AWLEN    (m8_awlen),
        .M8_AWSIZE   (m8_awsize),
        .M8_AWBURST  (m8_awburst),
        .M8_AWLOCK   (m8_awlock),
        .M8_AWCACHE  (m8_awcache),
        .M8_AWPROT   (m8_awprot),
        .M8_AWQOS    (m8_awqos),
        .M8_AWREGION (4'b0000),
        .M8_AWVALID  (m8_awvalid),
        .M8_AWREADY  (m8_awready),
        .M8_WDATA    (m8_wdata),
        .M8_WSTRB    (m8_wstrb),
        .M8_WLAST    (m8_wlast),
        .M8_WVALID   (m8_wvalid),
        .M8_WREADY   (m8_wready),
        .M8_BID      (m8_bid),
        .M8_BRESP    (m8_bresp),
        .M8_BVALID   (m8_bvalid),
        .M8_BREADY   (m8_bready),
        .M8_ARID     (m8_arid),
        .M8_ARADDR   (m8_araddr),
        .M8_ARLEN    (m8_arlen),
        .M8_ARSIZE   (m8_arsize),
        .M8_ARBURST  (m8_arburst),
        .M8_ARLOCK   (m8_arlock),
        .M8_ARCACHE  (m8_arcache),
        .M8_ARPROT   (m8_arprot),
        .M8_ARQOS    (m8_arqos),
        .M8_ARREGION (4'b0000),
        .M8_ARVALID  (m8_arvalid),
        .M8_ARREADY  (m8_arready),
        .M8_RID      (m8_rid),
        .M8_RDATA    (m8_rdata),
        .M8_RRESP    (m8_rresp),
        .M8_RLAST    (m8_rlast),
        .M8_RVALID   (m8_rvalid),
        .M8_RREADY   (m8_rready),
        
        // Slave 0
        .S0_AWID     (s0_awid),
        .S0_AWADDR   (s0_awaddr),
        .S0_AWLEN    (s0_awlen),
        .S0_AWSIZE   (s0_awsize),
        .S0_AWBURST  (s0_awburst),
        .S0_AWLOCK   (s0_awlock),
        .S0_AWCACHE  (s0_awcache),
        .S0_AWPROT   (s0_awprot),
        .S0_AWQOS    (s0_awqos),
        .S0_AWREGION (),  // Not connected
        .S0_AWVALID  (s0_awvalid),
        .S0_AWREADY  (s0_awready),
        .S0_WDATA    (s0_wdata),
        .S0_WSTRB    (s0_wstrb),
        .S0_WLAST    (s0_wlast),
        .S0_WVALID   (s0_wvalid),
        .S0_WREADY   (s0_wready),
        .S0_BID      (s0_bid),
        .S0_BRESP    (s0_bresp),
        .S0_BVALID   (s0_bvalid),
        .S0_BREADY   (s0_bready),
        .S0_ARID     (s0_arid),
        .S0_ARADDR   (s0_araddr),
        .S0_ARLEN    (s0_arlen),
        .S0_ARSIZE   (s0_arsize),
        .S0_ARBURST  (s0_arburst),
        .S0_ARLOCK   (s0_arlock),
        .S0_ARCACHE  (s0_arcache),
        .S0_ARPROT   (s0_arprot),
        .S0_ARQOS    (s0_arqos),
        .S0_ARREGION (),
        .S0_ARVALID  (s0_arvalid),
        .S0_ARREADY  (s0_arready),
        .S0_RID      (s0_rid),
        .S0_RDATA    (s0_rdata),
        .S0_RRESP    (s0_rresp),
        .S0_RLAST    (s0_rlast),
        .S0_RVALID   (s0_rvalid),
        .S0_RREADY   (s0_rready),
        
        // Slave 1
        .S1_AWID     (s1_awid),
        .S1_AWADDR   (s1_awaddr),
        .S1_AWLEN    (s1_awlen),
        .S1_AWSIZE   (s1_awsize),
        .S1_AWBURST  (s1_awburst),
        .S1_AWLOCK   (s1_awlock),
        .S1_AWCACHE  (s1_awcache),
        .S1_AWPROT   (s1_awprot),
        .S1_AWQOS    (s1_awqos),
        .S1_AWREGION (),
        .S1_AWVALID  (s1_awvalid),
        .S1_AWREADY  (s1_awready),
        .S1_WDATA    (s1_wdata),
        .S1_WSTRB    (s1_wstrb),
        .S1_WLAST    (s1_wlast),
        .S1_WVALID   (s1_wvalid),
        .S1_WREADY   (s1_wready),
        .S1_BID      (s1_bid),
        .S1_BRESP    (s1_bresp),
        .S1_BVALID   (s1_bvalid),
        .S1_BREADY   (s1_bready),
        .S1_ARID     (s1_arid),
        .S1_ARADDR   (s1_araddr),
        .S1_ARLEN    (s1_arlen),
        .S1_ARSIZE   (s1_arsize),
        .S1_ARBURST  (s1_arburst),
        .S1_ARLOCK   (s1_arlock),
        .S1_ARCACHE  (s1_arcache),
        .S1_ARPROT   (s1_arprot),
        .S1_ARQOS    (s1_arqos),
        .S1_ARREGION (),
        .S1_ARVALID  (s1_arvalid),
        .S1_ARREADY  (s1_arready),
        .S1_RID      (s1_rid),
        .S1_RDATA    (s1_rdata),
        .S1_RRESP    (s1_rresp),
        .S1_RLAST    (s1_rlast),
        .S1_RVALID   (s1_rvalid),
        .S1_RREADY   (s1_rready),
        
        // Slave 2
        .S2_AWID     (s2_awid),
        .S2_AWADDR   (s2_awaddr),
        .S2_AWLEN    (s2_awlen),
        .S2_AWSIZE   (s2_awsize),
        .S2_AWBURST  (s2_awburst),
        .S2_AWLOCK   (s2_awlock),
        .S2_AWCACHE  (s2_awcache),
        .S2_AWPROT   (s2_awprot),
        .S2_AWQOS    (s2_awqos),
        .S2_AWREGION (),
        .S2_AWVALID  (s2_awvalid),
        .S2_AWREADY  (s2_awready),
        .S2_WDATA    (s2_wdata),
        .S2_WSTRB    (s2_wstrb),
        .S2_WLAST    (s2_wlast),
        .S2_WVALID   (s2_wvalid),
        .S2_WREADY   (s2_wready),
        .S2_BID      (s2_bid),
        .S2_BRESP    (s2_bresp),
        .S2_BVALID   (s2_bvalid),
        .S2_BREADY   (s2_bready),
        .S2_ARID     (s2_arid),
        .S2_ARADDR   (s2_araddr),
        .S2_ARLEN    (s2_arlen),
        .S2_ARSIZE   (s2_arsize),
        .S2_ARBURST  (s2_arburst),
        .S2_ARLOCK   (s2_arlock),
        .S2_ARCACHE  (s2_arcache),
        .S2_ARPROT   (s2_arprot),
        .S2_ARQOS    (s2_arqos),
        .S2_ARREGION (),
        .S2_ARVALID  (s2_arvalid),
        .S2_ARREADY  (s2_arready),
        .S2_RID      (s2_rid),
        .S2_RDATA    (s2_rdata),
        .S2_RRESP    (s2_rresp),
        .S2_RLAST    (s2_rlast),
        .S2_RVALID   (s2_rvalid),
        .S2_RREADY   (s2_rready),
        
        // Slave 3
        .S3_AWID     (s3_awid),
        .S3_AWADDR   (s3_awaddr),
        .S3_AWLEN    (s3_awlen),
        .S3_AWSIZE   (s3_awsize),
        .S3_AWBURST  (s3_awburst),
        .S3_AWLOCK   (s3_awlock),
        .S3_AWCACHE  (s3_awcache),
        .S3_AWPROT   (s3_awprot),
        .S3_AWQOS    (s3_awqos),
        .S3_AWREGION (),
        .S3_AWVALID  (s3_awvalid),
        .S3_AWREADY  (s3_awready),
        .S3_WDATA    (s3_wdata),
        .S3_WSTRB    (s3_wstrb),
        .S3_WLAST    (s3_wlast),
        .S3_WVALID   (s3_wvalid),
        .S3_WREADY   (s3_wready),
        .S3_BID      (s3_bid),
        .S3_BRESP    (s3_bresp),
        .S3_BVALID   (s3_bvalid),
        .S3_BREADY   (s3_bready),
        .S3_ARID     (s3_arid),
        .S3_ARADDR   (s3_araddr),
        .S3_ARLEN    (s3_arlen),
        .S3_ARSIZE   (s3_arsize),
        .S3_ARBURST  (s3_arburst),
        .S3_ARLOCK   (s3_arlock),
        .S3_ARCACHE  (s3_arcache),
        .S3_ARPROT   (s3_arprot),
        .S3_ARQOS    (s3_arqos),
        .S3_ARREGION (),
        .S3_ARVALID  (s3_arvalid),
        .S3_ARREADY  (s3_arready),
        .S3_RID      (s3_rid),
        .S3_RDATA    (s3_rdata),
        .S3_RRESP    (s3_rresp),
        .S3_RLAST    (s3_rlast),
        .S3_RVALID   (s3_rvalid),
        .S3_RREADY   (s3_rready),
        
        // Slave 4
        .S4_AWID     (s4_awid),
        .S4_AWADDR   (s4_awaddr),
        .S4_AWLEN    (s4_awlen),
        .S4_AWSIZE   (s4_awsize),
        .S4_AWBURST  (s4_awburst),
        .S4_AWLOCK   (s4_awlock),
        .S4_AWCACHE  (s4_awcache),
        .S4_AWPROT   (s4_awprot),
        .S4_AWQOS    (s4_awqos),
        .S4_AWREGION (),
        .S4_AWVALID  (s4_awvalid),
        .S4_AWREADY  (s4_awready),
        .S4_WDATA    (s4_wdata),
        .S4_WSTRB    (s4_wstrb),
        .S4_WLAST    (s4_wlast),
        .S4_WVALID   (s4_wvalid),
        .S4_WREADY   (s4_wready),
        .S4_BID      (s4_bid),
        .S4_BRESP    (s4_bresp),
        .S4_BVALID   (s4_bvalid),
        .S4_BREADY   (s4_bready),
        .S4_ARID     (s4_arid),
        .S4_ARADDR   (s4_araddr),
        .S4_ARLEN    (s4_arlen),
        .S4_ARSIZE   (s4_arsize),
        .S4_ARBURST  (s4_arburst),
        .S4_ARLOCK   (s4_arlock),
        .S4_ARCACHE  (s4_arcache),
        .S4_ARPROT   (s4_arprot),
        .S4_ARQOS    (s4_arqos),
        .S4_ARREGION (),
        .S4_ARVALID  (s4_arvalid),
        .S4_ARREADY  (s4_arready),
        .S4_RID      (s4_rid),
        .S4_RDATA    (s4_rdata),
        .S4_RRESP    (s4_rresp),
        .S4_RLAST    (s4_rlast),
        .S4_RVALID   (s4_rvalid),
        .S4_RREADY   (s4_rready),
        
        // Slave 5
        .S5_AWID     (s5_awid),
        .S5_AWADDR   (s5_awaddr),
        .S5_AWLEN    (s5_awlen),
        .S5_AWSIZE   (s5_awsize),
        .S5_AWBURST  (s5_awburst),
        .S5_AWLOCK   (s5_awlock),
        .S5_AWCACHE  (s5_awcache),
        .S5_AWPROT   (s5_awprot),
        .S5_AWQOS    (s5_awqos),
        .S5_AWREGION (),
        .S5_AWVALID  (s5_awvalid),
        .S5_AWREADY  (s5_awready),
        .S5_WDATA    (s5_wdata),
        .S5_WSTRB    (s5_wstrb),
        .S5_WLAST    (s5_wlast),
        .S5_WVALID   (s5_wvalid),
        .S5_WREADY   (s5_wready),
        .S5_BID      (s5_bid),
        .S5_BRESP    (s5_bresp),
        .S5_BVALID   (s5_bvalid),
        .S5_BREADY   (s5_bready),
        .S5_ARID     (s5_arid),
        .S5_ARADDR   (s5_araddr),
        .S5_ARLEN    (s5_arlen),
        .S5_ARSIZE   (s5_arsize),
        .S5_ARBURST  (s5_arburst),
        .S5_ARLOCK   (s5_arlock),
        .S5_ARCACHE  (s5_arcache),
        .S5_ARPROT   (s5_arprot),
        .S5_ARQOS    (s5_arqos),
        .S5_ARREGION (),
        .S5_ARVALID  (s5_arvalid),
        .S5_ARREADY  (s5_arready),
        .S5_RID      (s5_rid),
        .S5_RDATA    (s5_rdata),
        .S5_RRESP    (s5_rresp),
        .S5_RLAST    (s5_rlast),
        .S5_RVALID   (s5_rvalid),
        .S5_RREADY   (s5_rready),
        
        // Slave 6
        .S6_AWID     (s6_awid),
        .S6_AWADDR   (s6_awaddr),
        .S6_AWLEN    (s6_awlen),
        .S6_AWSIZE   (s6_awsize),
        .S6_AWBURST  (s6_awburst),
        .S6_AWLOCK   (s6_awlock),
        .S6_AWCACHE  (s6_awcache),
        .S6_AWPROT   (s6_awprot),
        .S6_AWQOS    (s6_awqos),
        .S6_AWREGION (),
        .S6_AWVALID  (s6_awvalid),
        .S6_AWREADY  (s6_awready),
        .S6_WDATA    (s6_wdata),
        .S6_WSTRB    (s6_wstrb),
        .S6_WLAST    (s6_wlast),
        .S6_WVALID   (s6_wvalid),
        .S6_WREADY   (s6_wready),
        .S6_BID      (s6_bid),
        .S6_BRESP    (s6_bresp),
        .S6_BVALID   (s6_bvalid),
        .S6_BREADY   (s6_bready),
        .S6_ARID     (s6_arid),
        .S6_ARADDR   (s6_araddr),
        .S6_ARLEN    (s6_arlen),
        .S6_ARSIZE   (s6_arsize),
        .S6_ARBURST  (s6_arburst),
        .S6_ARLOCK   (s6_arlock),
        .S6_ARCACHE  (s6_arcache),
        .S6_ARPROT   (s6_arprot),
        .S6_ARQOS    (s6_arqos),
        .S6_ARREGION (),
        .S6_ARVALID  (s6_arvalid),
        .S6_ARREADY  (s6_arready),
        .S6_RID      (s6_rid),
        .S6_RDATA    (s6_rdata),
        .S6_RRESP    (s6_rresp),
        .S6_RLAST    (s6_rlast),
        .S6_RVALID   (s6_rvalid),
        .S6_RREADY   (s6_rready),
        
        // Slave 7
        .S7_AWID     (s7_awid),
        .S7_AWADDR   (s7_awaddr),
        .S7_AWLEN    (s7_awlen),
        .S7_AWSIZE   (s7_awsize),
        .S7_AWBURST  (s7_awburst),
        .S7_AWLOCK   (s7_awlock),
        .S7_AWCACHE  (s7_awcache),
        .S7_AWPROT   (s7_awprot),
        .S7_AWQOS    (s7_awqos),
        .S7_AWREGION (),
        .S7_AWVALID  (s7_awvalid),
        .S7_AWREADY  (s7_awready),
        .S7_WDATA    (s7_wdata),
        .S7_WSTRB    (s7_wstrb),
        .S7_WLAST    (s7_wlast),
        .S7_WVALID   (s7_wvalid),
        .S7_WREADY   (s7_wready),
        .S7_BID      (s7_bid),
        .S7_BRESP    (s7_bresp),
        .S7_BVALID   (s7_bvalid),
        .S7_BREADY   (s7_bready),
        .S7_ARID     (s7_arid),
        .S7_ARADDR   (s7_araddr),
        .S7_ARLEN    (s7_arlen),
        .S7_ARSIZE   (s7_arsize),
        .S7_ARBURST  (s7_arburst),
        .S7_ARLOCK   (s7_arlock),
        .S7_ARCACHE  (s7_arcache),
        .S7_ARPROT   (s7_arprot),
        .S7_ARQOS    (s7_arqos),
        .S7_ARREGION (),
        .S7_ARVALID  (s7_arvalid),
        .S7_ARREADY  (s7_arready),
        .S7_RID      (s7_rid),
        .S7_RDATA    (s7_rdata),
        .S7_RRESP    (s7_rresp),
        .S7_RLAST    (s7_rlast),
        .S7_RVALID   (s7_rvalid),
        .S7_RREADY   (s7_rready),
        
        // Slave 8
        .S8_AWID     (s8_awid),
        .S8_AWADDR   (s8_awaddr),
        .S8_AWLEN    (s8_awlen),
        .S8_AWSIZE   (s8_awsize),
        .S8_AWBURST  (s8_awburst),
        .S8_AWLOCK   (s8_awlock),
        .S8_AWCACHE  (s8_awcache),
        .S8_AWPROT   (s8_awprot),
        .S8_AWQOS    (s8_awqos),
        .S8_AWREGION (),
        .S8_AWVALID  (s8_awvalid),
        .S8_AWREADY  (s8_awready),
        .S8_WDATA    (s8_wdata),
        .S8_WSTRB    (s8_wstrb),
        .S8_WLAST    (s8_wlast),
        .S8_WVALID   (s8_wvalid),
        .S8_WREADY   (s8_wready),
        .S8_BID      (s8_bid),
        .S8_BRESP    (s8_bresp),
        .S8_BVALID   (s8_bvalid),
        .S8_BREADY   (s8_bready),
        .S8_ARID     (s8_arid),
        .S8_ARADDR   (s8_araddr),
        .S8_ARLEN    (s8_arlen),
        .S8_ARSIZE   (s8_arsize),
        .S8_ARBURST  (s8_arburst),
        .S8_ARLOCK   (s8_arlock),
        .S8_ARCACHE  (s8_arcache),
        .S8_ARPROT   (s8_arprot),
        .S8_ARQOS    (s8_arqos),
        .S8_ARREGION (),
        .S8_ARVALID  (s8_arvalid),
        .S8_ARREADY  (s8_arready),
        .S8_RID      (s8_rid),
        .S8_RDATA    (s8_rdata),
        .S8_RRESP    (s8_rresp),
        .S8_RLAST    (s8_rlast),
        .S8_RVALID   (s8_rvalid),
        .S8_RREADY   (s8_rready)
    );

endmodule