// Master wire declarations for Masters 1-14
// This file is included in dut_wrapper_real_rtl.sv

// Master 1
wire [RTL_ID_WIDTH-1:0]     m1_awid;
wire [ADDR_WIDTH-1:0]       m1_awaddr;
wire [7:0]                  m1_awlen;
wire [2:0]                  m1_awsize;
wire [1:0]                  m1_awburst;
wire                        m1_awlock;
wire [3:0]                  m1_awcache;
wire [2:0]                  m1_awprot;
wire [3:0]                  m1_awqos;
wire                        m1_awvalid;
wire                        m1_awready;
wire [DATA_WIDTH-1:0]       m1_wdata;
wire [DATA_WIDTH/8-1:0]     m1_wstrb;
wire                        m1_wlast;
wire                        m1_wvalid;
wire                        m1_wready;
wire [RTL_ID_WIDTH-1:0]     m1_bid;
wire [1:0]                  m1_bresp;
wire                        m1_bvalid;
wire                        m1_bready;
wire [RTL_ID_WIDTH-1:0]     m1_arid;
wire [ADDR_WIDTH-1:0]       m1_araddr;
wire [7:0]                  m1_arlen;
wire [2:0]                  m1_arsize;
wire [1:0]                  m1_arburst;
wire                        m1_arlock;
wire [3:0]                  m1_arcache;
wire [2:0]                  m1_arprot;
wire [3:0]                  m1_arqos;
wire                        m1_arvalid;
wire                        m1_arready;
wire [RTL_ID_WIDTH-1:0]     m1_rid;
wire [DATA_WIDTH-1:0]       m1_rdata;
wire [1:0]                  m1_rresp;
wire                        m1_rlast;
wire                        m1_rvalid;
wire                        m1_rready;

// Master 2
wire [RTL_ID_WIDTH-1:0]     m2_awid;
wire [ADDR_WIDTH-1:0]       m2_awaddr;
wire [7:0]                  m2_awlen;
wire [2:0]                  m2_awsize;
wire [1:0]                  m2_awburst;
wire                        m2_awlock;
wire [3:0]                  m2_awcache;
wire [2:0]                  m2_awprot;
wire [3:0]                  m2_awqos;
wire                        m2_awvalid;
wire                        m2_awready;
wire [DATA_WIDTH-1:0]       m2_wdata;
wire [DATA_WIDTH/8-1:0]     m2_wstrb;
wire                        m2_wlast;
wire                        m2_wvalid;
wire                        m2_wready;
wire [RTL_ID_WIDTH-1:0]     m2_bid;
wire [1:0]                  m2_bresp;
wire                        m2_bvalid;
wire                        m2_bready;
wire [RTL_ID_WIDTH-1:0]     m2_arid;
wire [ADDR_WIDTH-1:0]       m2_araddr;
wire [7:0]                  m2_arlen;
wire [2:0]                  m2_arsize;
wire [1:0]                  m2_arburst;
wire                        m2_arlock;
wire [3:0]                  m2_arcache;
wire [2:0]                  m2_arprot;
wire [3:0]                  m2_arqos;
wire                        m2_arvalid;
wire                        m2_arready;
wire [RTL_ID_WIDTH-1:0]     m2_rid;
wire [DATA_WIDTH-1:0]       m2_rdata;
wire [1:0]                  m2_rresp;
wire                        m2_rlast;
wire                        m2_rvalid;
wire                        m2_rready;

// Master 3
wire [RTL_ID_WIDTH-1:0]     m3_awid;
wire [ADDR_WIDTH-1:0]       m3_awaddr;
wire [7:0]                  m3_awlen;
wire [2:0]                  m3_awsize;
wire [1:0]                  m3_awburst;
wire                        m3_awlock;
wire [3:0]                  m3_awcache;
wire [2:0]                  m3_awprot;
wire [3:0]                  m3_awqos;
wire                        m3_awvalid;
wire                        m3_awready;
wire [DATA_WIDTH-1:0]       m3_wdata;
wire [DATA_WIDTH/8-1:0]     m3_wstrb;
wire                        m3_wlast;
wire                        m3_wvalid;
wire                        m3_wready;
wire [RTL_ID_WIDTH-1:0]     m3_bid;
wire [1:0]                  m3_bresp;
wire                        m3_bvalid;
wire                        m3_bready;
wire [RTL_ID_WIDTH-1:0]     m3_arid;
wire [ADDR_WIDTH-1:0]       m3_araddr;
wire [7:0]                  m3_arlen;
wire [2:0]                  m3_arsize;
wire [1:0]                  m3_arburst;
wire                        m3_arlock;
wire [3:0]                  m3_arcache;
wire [2:0]                  m3_arprot;
wire [3:0]                  m3_arqos;
wire                        m3_arvalid;
wire                        m3_arready;
wire [RTL_ID_WIDTH-1:0]     m3_rid;
wire [DATA_WIDTH-1:0]       m3_rdata;
wire [1:0]                  m3_rresp;
wire                        m3_rlast;
wire                        m3_rvalid;
wire                        m3_rready;

// Master 4
wire [RTL_ID_WIDTH-1:0]     m4_awid;
wire [ADDR_WIDTH-1:0]       m4_awaddr;
wire [7:0]                  m4_awlen;
wire [2:0]                  m4_awsize;
wire [1:0]                  m4_awburst;
wire                        m4_awlock;
wire [3:0]                  m4_awcache;
wire [2:0]                  m4_awprot;
wire [3:0]                  m4_awqos;
wire                        m4_awvalid;
wire                        m4_awready;
wire [DATA_WIDTH-1:0]       m4_wdata;
wire [DATA_WIDTH/8-1:0]     m4_wstrb;
wire                        m4_wlast;
wire                        m4_wvalid;
wire                        m4_wready;
wire [RTL_ID_WIDTH-1:0]     m4_bid;
wire [1:0]                  m4_bresp;
wire                        m4_bvalid;
wire                        m4_bready;
wire [RTL_ID_WIDTH-1:0]     m4_arid;
wire [ADDR_WIDTH-1:0]       m4_araddr;
wire [7:0]                  m4_arlen;
wire [2:0]                  m4_arsize;
wire [1:0]                  m4_arburst;
wire                        m4_arlock;
wire [3:0]                  m4_arcache;
wire [2:0]                  m4_arprot;
wire [3:0]                  m4_arqos;
wire                        m4_arvalid;
wire                        m4_arready;
wire [RTL_ID_WIDTH-1:0]     m4_rid;
wire [DATA_WIDTH-1:0]       m4_rdata;
wire [1:0]                  m4_rresp;
wire                        m4_rlast;
wire                        m4_rvalid;
wire                        m4_rready;

// Master 5
wire [RTL_ID_WIDTH-1:0]     m5_awid;
wire [ADDR_WIDTH-1:0]       m5_awaddr;
wire [7:0]                  m5_awlen;
wire [2:0]                  m5_awsize;
wire [1:0]                  m5_awburst;
wire                        m5_awlock;
wire [3:0]                  m5_awcache;
wire [2:0]                  m5_awprot;
wire [3:0]                  m5_awqos;
wire                        m5_awvalid;
wire                        m5_awready;
wire [DATA_WIDTH-1:0]       m5_wdata;
wire [DATA_WIDTH/8-1:0]     m5_wstrb;
wire                        m5_wlast;
wire                        m5_wvalid;
wire                        m5_wready;
wire [RTL_ID_WIDTH-1:0]     m5_bid;
wire [1:0]                  m5_bresp;
wire                        m5_bvalid;
wire                        m5_bready;
wire [RTL_ID_WIDTH-1:0]     m5_arid;
wire [ADDR_WIDTH-1:0]       m5_araddr;
wire [7:0]                  m5_arlen;
wire [2:0]                  m5_arsize;
wire [1:0]                  m5_arburst;
wire                        m5_arlock;
wire [3:0]                  m5_arcache;
wire [2:0]                  m5_arprot;
wire [3:0]                  m5_arqos;
wire                        m5_arvalid;
wire                        m5_arready;
wire [RTL_ID_WIDTH-1:0]     m5_rid;
wire [DATA_WIDTH-1:0]       m5_rdata;
wire [1:0]                  m5_rresp;
wire                        m5_rlast;
wire                        m5_rvalid;
wire                        m5_rready;

// Master 6
wire [RTL_ID_WIDTH-1:0]     m6_awid;
wire [ADDR_WIDTH-1:0]       m6_awaddr;
wire [7:0]                  m6_awlen;
wire [2:0]                  m6_awsize;
wire [1:0]                  m6_awburst;
wire                        m6_awlock;
wire [3:0]                  m6_awcache;
wire [2:0]                  m6_awprot;
wire [3:0]                  m6_awqos;
wire                        m6_awvalid;
wire                        m6_awready;
wire [DATA_WIDTH-1:0]       m6_wdata;
wire [DATA_WIDTH/8-1:0]     m6_wstrb;
wire                        m6_wlast;
wire                        m6_wvalid;
wire                        m6_wready;
wire [RTL_ID_WIDTH-1:0]     m6_bid;
wire [1:0]                  m6_bresp;
wire                        m6_bvalid;
wire                        m6_bready;
wire [RTL_ID_WIDTH-1:0]     m6_arid;
wire [ADDR_WIDTH-1:0]       m6_araddr;
wire [7:0]                  m6_arlen;
wire [2:0]                  m6_arsize;
wire [1:0]                  m6_arburst;
wire                        m6_arlock;
wire [3:0]                  m6_arcache;
wire [2:0]                  m6_arprot;
wire [3:0]                  m6_arqos;
wire                        m6_arvalid;
wire                        m6_arready;
wire [RTL_ID_WIDTH-1:0]     m6_rid;
wire [DATA_WIDTH-1:0]       m6_rdata;
wire [1:0]                  m6_rresp;
wire                        m6_rlast;
wire                        m6_rvalid;
wire                        m6_rready;

// Master 7
wire [RTL_ID_WIDTH-1:0]     m7_awid;
wire [ADDR_WIDTH-1:0]       m7_awaddr;
wire [7:0]                  m7_awlen;
wire [2:0]                  m7_awsize;
wire [1:0]                  m7_awburst;
wire                        m7_awlock;
wire [3:0]                  m7_awcache;
wire [2:0]                  m7_awprot;
wire [3:0]                  m7_awqos;
wire                        m7_awvalid;
wire                        m7_awready;
wire [DATA_WIDTH-1:0]       m7_wdata;
wire [DATA_WIDTH/8-1:0]     m7_wstrb;
wire                        m7_wlast;
wire                        m7_wvalid;
wire                        m7_wready;
wire [RTL_ID_WIDTH-1:0]     m7_bid;
wire [1:0]                  m7_bresp;
wire                        m7_bvalid;
wire                        m7_bready;
wire [RTL_ID_WIDTH-1:0]     m7_arid;
wire [ADDR_WIDTH-1:0]       m7_araddr;
wire [7:0]                  m7_arlen;
wire [2:0]                  m7_arsize;
wire [1:0]                  m7_arburst;
wire                        m7_arlock;
wire [3:0]                  m7_arcache;
wire [2:0]                  m7_arprot;
wire [3:0]                  m7_arqos;
wire                        m7_arvalid;
wire                        m7_arready;
wire [RTL_ID_WIDTH-1:0]     m7_rid;
wire [DATA_WIDTH-1:0]       m7_rdata;
wire [1:0]                  m7_rresp;
wire                        m7_rlast;
wire                        m7_rvalid;
wire                        m7_rready;

// Master 8
wire [RTL_ID_WIDTH-1:0]     m8_awid;
wire [ADDR_WIDTH-1:0]       m8_awaddr;
wire [7:0]                  m8_awlen;
wire [2:0]                  m8_awsize;
wire [1:0]                  m8_awburst;
wire                        m8_awlock;
wire [3:0]                  m8_awcache;
wire [2:0]                  m8_awprot;
wire [3:0]                  m8_awqos;
wire                        m8_awvalid;
wire                        m8_awready;
wire [DATA_WIDTH-1:0]       m8_wdata;
wire [DATA_WIDTH/8-1:0]     m8_wstrb;
wire                        m8_wlast;
wire                        m8_wvalid;
wire                        m8_wready;
wire [RTL_ID_WIDTH-1:0]     m8_bid;
wire [1:0]                  m8_bresp;
wire                        m8_bvalid;
wire                        m8_bready;
wire [RTL_ID_WIDTH-1:0]     m8_arid;
wire [ADDR_WIDTH-1:0]       m8_araddr;
wire [7:0]                  m8_arlen;
wire [2:0]                  m8_arsize;
wire [1:0]                  m8_arburst;
wire                        m8_arlock;
wire [3:0]                  m8_arcache;
wire [2:0]                  m8_arprot;
wire [3:0]                  m8_arqos;
wire                        m8_arvalid;
wire                        m8_arready;
wire [RTL_ID_WIDTH-1:0]     m8_rid;
wire [DATA_WIDTH-1:0]       m8_rdata;
wire [1:0]                  m8_rresp;
wire                        m8_rlast;
wire                        m8_rvalid;
wire                        m8_rready;

// Master 9
wire [RTL_ID_WIDTH-1:0]     m9_awid;
wire [ADDR_WIDTH-1:0]       m9_awaddr;
wire [7:0]                  m9_awlen;
wire [2:0]                  m9_awsize;
wire [1:0]                  m9_awburst;
wire                        m9_awlock;
wire [3:0]                  m9_awcache;
wire [2:0]                  m9_awprot;
wire [3:0]                  m9_awqos;
wire                        m9_awvalid;
wire                        m9_awready;
wire [DATA_WIDTH-1:0]       m9_wdata;
wire [DATA_WIDTH/8-1:0]     m9_wstrb;
wire                        m9_wlast;
wire                        m9_wvalid;
wire                        m9_wready;
wire [RTL_ID_WIDTH-1:0]     m9_bid;
wire [1:0]                  m9_bresp;
wire                        m9_bvalid;
wire                        m9_bready;
wire [RTL_ID_WIDTH-1:0]     m9_arid;
wire [ADDR_WIDTH-1:0]       m9_araddr;
wire [7:0]                  m9_arlen;
wire [2:0]                  m9_arsize;
wire [1:0]                  m9_arburst;
wire                        m9_arlock;
wire [3:0]                  m9_arcache;
wire [2:0]                  m9_arprot;
wire [3:0]                  m9_arqos;
wire                        m9_arvalid;
wire                        m9_arready;
wire [RTL_ID_WIDTH-1:0]     m9_rid;
wire [DATA_WIDTH-1:0]       m9_rdata;
wire [1:0]                  m9_rresp;
wire                        m9_rlast;
wire                        m9_rvalid;
wire                        m9_rready;

// Master 10
wire [RTL_ID_WIDTH-1:0]     m10_awid;
wire [ADDR_WIDTH-1:0]       m10_awaddr;
wire [7:0]                  m10_awlen;
wire [2:0]                  m10_awsize;
wire [1:0]                  m10_awburst;
wire                        m10_awlock;
wire [3:0]                  m10_awcache;
wire [2:0]                  m10_awprot;
wire [3:0]                  m10_awqos;
wire                        m10_awvalid;
wire                        m10_awready;
wire [DATA_WIDTH-1:0]       m10_wdata;
wire [DATA_WIDTH/8-1:0]     m10_wstrb;
wire                        m10_wlast;
wire                        m10_wvalid;
wire                        m10_wready;
wire [RTL_ID_WIDTH-1:0]     m10_bid;
wire [1:0]                  m10_bresp;
wire                        m10_bvalid;
wire                        m10_bready;
wire [RTL_ID_WIDTH-1:0]     m10_arid;
wire [ADDR_WIDTH-1:0]       m10_araddr;
wire [7:0]                  m10_arlen;
wire [2:0]                  m10_arsize;
wire [1:0]                  m10_arburst;
wire                        m10_arlock;
wire [3:0]                  m10_arcache;
wire [2:0]                  m10_arprot;
wire [3:0]                  m10_arqos;
wire                        m10_arvalid;
wire                        m10_arready;
wire [RTL_ID_WIDTH-1:0]     m10_rid;
wire [DATA_WIDTH-1:0]       m10_rdata;
wire [1:0]                  m10_rresp;
wire                        m10_rlast;
wire                        m10_rvalid;
wire                        m10_rready;

// Master 11
wire [RTL_ID_WIDTH-1:0]     m11_awid;
wire [ADDR_WIDTH-1:0]       m11_awaddr;
wire [7:0]                  m11_awlen;
wire [2:0]                  m11_awsize;
wire [1:0]                  m11_awburst;
wire                        m11_awlock;
wire [3:0]                  m11_awcache;
wire [2:0]                  m11_awprot;
wire [3:0]                  m11_awqos;
wire                        m11_awvalid;
wire                        m11_awready;
wire [DATA_WIDTH-1:0]       m11_wdata;
wire [DATA_WIDTH/8-1:0]     m11_wstrb;
wire                        m11_wlast;
wire                        m11_wvalid;
wire                        m11_wready;
wire [RTL_ID_WIDTH-1:0]     m11_bid;
wire [1:0]                  m11_bresp;
wire                        m11_bvalid;
wire                        m11_bready;
wire [RTL_ID_WIDTH-1:0]     m11_arid;
wire [ADDR_WIDTH-1:0]       m11_araddr;
wire [7:0]                  m11_arlen;
wire [2:0]                  m11_arsize;
wire [1:0]                  m11_arburst;
wire                        m11_arlock;
wire [3:0]                  m11_arcache;
wire [2:0]                  m11_arprot;
wire [3:0]                  m11_arqos;
wire                        m11_arvalid;
wire                        m11_arready;
wire [RTL_ID_WIDTH-1:0]     m11_rid;
wire [DATA_WIDTH-1:0]       m11_rdata;
wire [1:0]                  m11_rresp;
wire                        m11_rlast;
wire                        m11_rvalid;
wire                        m11_rready;

// Master 12
wire [RTL_ID_WIDTH-1:0]     m12_awid;
wire [ADDR_WIDTH-1:0]       m12_awaddr;
wire [7:0]                  m12_awlen;
wire [2:0]                  m12_awsize;
wire [1:0]                  m12_awburst;
wire                        m12_awlock;
wire [3:0]                  m12_awcache;
wire [2:0]                  m12_awprot;
wire [3:0]                  m12_awqos;
wire                        m12_awvalid;
wire                        m12_awready;
wire [DATA_WIDTH-1:0]       m12_wdata;
wire [DATA_WIDTH/8-1:0]     m12_wstrb;
wire                        m12_wlast;
wire                        m12_wvalid;
wire                        m12_wready;
wire [RTL_ID_WIDTH-1:0]     m12_bid;
wire [1:0]                  m12_bresp;
wire                        m12_bvalid;
wire                        m12_bready;
wire [RTL_ID_WIDTH-1:0]     m12_arid;
wire [ADDR_WIDTH-1:0]       m12_araddr;
wire [7:0]                  m12_arlen;
wire [2:0]                  m12_arsize;
wire [1:0]                  m12_arburst;
wire                        m12_arlock;
wire [3:0]                  m12_arcache;
wire [2:0]                  m12_arprot;
wire [3:0]                  m12_arqos;
wire                        m12_arvalid;
wire                        m12_arready;
wire [RTL_ID_WIDTH-1:0]     m12_rid;
wire [DATA_WIDTH-1:0]       m12_rdata;
wire [1:0]                  m12_rresp;
wire                        m12_rlast;
wire                        m12_rvalid;
wire                        m12_rready;

// Master 13
wire [RTL_ID_WIDTH-1:0]     m13_awid;
wire [ADDR_WIDTH-1:0]       m13_awaddr;
wire [7:0]                  m13_awlen;
wire [2:0]                  m13_awsize;
wire [1:0]                  m13_awburst;
wire                        m13_awlock;
wire [3:0]                  m13_awcache;
wire [2:0]                  m13_awprot;
wire [3:0]                  m13_awqos;
wire                        m13_awvalid;
wire                        m13_awready;
wire [DATA_WIDTH-1:0]       m13_wdata;
wire [DATA_WIDTH/8-1:0]     m13_wstrb;
wire                        m13_wlast;
wire                        m13_wvalid;
wire                        m13_wready;
wire [RTL_ID_WIDTH-1:0]     m13_bid;
wire [1:0]                  m13_bresp;
wire                        m13_bvalid;
wire                        m13_bready;
wire [RTL_ID_WIDTH-1:0]     m13_arid;
wire [ADDR_WIDTH-1:0]       m13_araddr;
wire [7:0]                  m13_arlen;
wire [2:0]                  m13_arsize;
wire [1:0]                  m13_arburst;
wire                        m13_arlock;
wire [3:0]                  m13_arcache;
wire [2:0]                  m13_arprot;
wire [3:0]                  m13_arqos;
wire                        m13_arvalid;
wire                        m13_arready;
wire [RTL_ID_WIDTH-1:0]     m13_rid;
wire [DATA_WIDTH-1:0]       m13_rdata;
wire [1:0]                  m13_rresp;
wire                        m13_rlast;
wire                        m13_rvalid;
wire                        m13_rready;

// Master 14
wire [RTL_ID_WIDTH-1:0]     m14_awid;
wire [ADDR_WIDTH-1:0]       m14_awaddr;
wire [7:0]                  m14_awlen;
wire [2:0]                  m14_awsize;
wire [1:0]                  m14_awburst;
wire                        m14_awlock;
wire [3:0]                  m14_awcache;
wire [2:0]                  m14_awprot;
wire [3:0]                  m14_awqos;
wire                        m14_awvalid;
wire                        m14_awready;
wire [DATA_WIDTH-1:0]       m14_wdata;
wire [DATA_WIDTH/8-1:0]     m14_wstrb;
wire                        m14_wlast;
wire                        m14_wvalid;
wire                        m14_wready;
wire [RTL_ID_WIDTH-1:0]     m14_bid;
wire [1:0]                  m14_bresp;
wire                        m14_bvalid;
wire                        m14_bready;
wire [RTL_ID_WIDTH-1:0]     m14_arid;
wire [ADDR_WIDTH-1:0]       m14_araddr;
wire [7:0]                  m14_arlen;
wire [2:0]                  m14_arsize;
wire [1:0]                  m14_arburst;
wire                        m14_arlock;
wire [3:0]                  m14_arcache;
wire [2:0]                  m14_arprot;
wire [3:0]                  m14_arqos;
wire                        m14_arvalid;
wire                        m14_arready;
wire [RTL_ID_WIDTH-1:0]     m14_rid;
wire [DATA_WIDTH-1:0]       m14_rdata;
wire [1:0]                  m14_rresp;
wire                        m14_rlast;
wire                        m14_rvalid;
wire                        m14_rready;